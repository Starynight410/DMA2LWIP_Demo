`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Jo0GTP48lurGV9QI1c62RTUP1YVEamMz1VZFzIOsgfj+B/Me/Uz/+TNhvOgX00Boh3rVDWY3miWC
6dvD9WUK3Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LQaetkHlTEQ/O2QuW4ImDf/K0WBzrX60Y2eOh0Fzlit7V6+gYpu/pdjpcV2iUJ0OSkPSJI+Mhtnw
My00nmvcw7hr27JQMftgpSq2KJTPiuvMTKQgaTjH7G11dDQzZg5OIfVuhiEdrvLjBL6ODFpLjnot
+wtza061w0h0SULGF8g=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e7yz9u7SkKHpUf45ToebPKpSB+7SYjKyIPDWMVo4RpE1fApRY5i+m6AdkyczFN3egPL9yuxMUBQi
B3fcWe1KL481lABpqgSqODHUHO2V3VOpcYtVbs+ITdbbKzYLqgggxX2OFaFxfaKpm8KQDKkYwb5s
hDH0bmxkegiSbK8/6cCO7THsM2QEi5MCtiINLnSFKZxzW2n5D4XuM/reG5kcwrmcvNmgwL09iDms
zsLNFk+KlTwGLQ+sjNp4XMp3wRVy8au+yG/ZaAjv1SaonTr0s0Ktoq7kpKzzK8Vdx3gxl98oC7lG
qI6lKENHTJsj2Et1sJqARwUVTfXhIwUnx7z+eQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YUgiCLqe/j/NhPlORdPixdVwbLBtEL3BY6gCgf7tGi15P5FTCSoEIKV1fMOt5n55kUiULz6ixyOx
w6KSNkCTxNK1tRyjWlYPNwh+30X1DX2lqxQedujI8dEfW4TThaFzjbr5VzZ5Xx3QklpDtemVWlfc
v+85sRR7dpK2+yz7JHTpwsBUmUIz/yQuKTPH3TXkcTEtK3SDtuMd9W57I7EJRQs/QWb0HRC1gqri
b73Bznz/ITOHvk6hyVhz2IcLVxpPIWw2SPni76CtRBGxpvEkYBsB4Tb29iojsozDmdeCBCdMwy/R
z6g42MtTw4HdwvXecIHU1Ps+g//YLogOmAG9jA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
m7rYtXUavsevrUPbAA9ErlXCOGGk4fAoeRrucNOvvuTkTuigciZtMDGFuNCCP84AUenq7yf+knfr
YxGJdpaWbSksXpHqc2OaU9JxiGbOYXsVLB6aaIcsBViJ1Iu9Y3dsxqVRuEf/+KOaUoj9MgYpzlBd
dGJCSN02BKWDuiELCvkTzxH0HkaQw6L4Fs4eaqtvZO6JC37ps+GYsLvCsUVOUrxP3ZXffR/5rO+/
r+Y7T74S//4yP9CGXNTnVBNea7FKmyEzggzbDLVXfwg7DC9jqBdVLhJdArtJhH0AWfbyCLDAfF69
TIFn/nOkcwqHGmFmfhdLuMOHq1GabkUC03gqCw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WkzTVLle3kbJDg7jpvQ16rMwFjgKsN6s5VraGMgY5PuWLmuM4CseW8hGJcsf4WjZloefR1XKRkv+
EV0MnXlsj7dM99Z1mYpSYEt+FSSlVw8ZrTFDfAXM2tVaQ6tHWq2thbcjDszMiCZNwxeaVwffojNF
dPRWtPW7gJ6hRMZJ1oE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nB0LvvHetoBgxBsMSEPN44HAKokSVtsq+whVeE4wsASFbqJ8K82xM3hbmxu6ZDYkwRj1/AOA3HVk
G4ilfKGLy/G7TDbQDfRO+5Y01cbhrcP/GMxbBzv8olyMaD/JTd0uTncjO8AIV8tUE18Kj9ZhfRCb
zatytXSeRs9JZ1gbnMMyuS9DWHly6IquSzk4ICOoWWjyjXwHRFPGPkYHKeAKIXuBgNn5YIUb73Bg
ZfSxBEDnDG4lR9r5BsXVWXPmkRPzzmalgCEOM4dNamRFXJG6Z063apEzsaFADjlPswBxcO39daPt
PO0nWMUFnDtLtq5NhL5JcY8vaGgEnfVUj0929g==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kx2/4FUG+WgpOeMb3Rbb/cih1lc163wBQ4vKkckklmR615Brrk0uvh47GWx5YPIQIJ1dUYGfGof0
suWssmlsLprBF4iyZ0oJN+doxvhmSoNuyqNtF4sOBh2mA2fEVAiuuRzdRQMw/lsxuNxU5tTeu4Hq
m6fseqlUS4i/DqAjB6NT+vlMZPYsrIaV5xH4A+ZthsSp/Yv1VhT2z1Yf0I1zXIDSJLePBat4WiXu
ztJa66W8SRYkuIFjEUecZElA0JE2MfS3tIGvepvw+Jw2NqcpRNOyHazWtDF1qGPoplQ2+iAwhvFE
swC4IvCafgzOO12FbZwI5Wi1IC0+7hrnR+7e/A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
8GvLC41uBcFwr5Ki5OvQAwh2MwnGKfuE0FkJhaohC6KDT4SH9pKcwnvFqbHTm7H+kxpfjlg3NYlo
R8dPW4XArskiR6Di2uUoB/KHQZgA9Q3EtCXwkVLVQYGosg4UrfQHBMy+RfyZEy92HGHNUxOrd6ID
xlrs459kSET88zsv2Ay7STCfvwufPDyyNcSCFsXWfT6R+72IX/rABNjwcgY/Oo0uWWEoVWlXEQaa
8tsY+Au92TptzKnO/T9WpKKqtfqmJcy+zwcxj1cenRTwtg+v1Ibpj9LPeXj5eqUtN77hR1dtw/ll
2bu3pdhGvi6UQyNubOIk9DkNm/GtOEWxyQo2XjnAzjJi/4t2NamtqBVSlKWB1uUoZau/Q/UeaJRg
nSnoclzhI5OXUklMJozygiF5hTWRQtLqkcVQ766JZKSayNe47xZ49JhFkFQHTS2xrMp7AS4P4Wjq
IVjbtY4RJzTrBT2+tLAsWNrNENo85bxXeIVKRpyVDtaXjoFHcl6mGHuXofIj4Sn62ujjfEJhmP3V
5zfnW2ryuYrTb3JqoYNZn6dDAZs/WwTI4F5RG9gCYbLIJwkYpH6fH/gDFbiXcIYXk3ldWDcEpZse
pF0AQMwU6TsdC6FfZyD4CQpPhSpHGIQeRJlS4+ADHW2nT43A9XuUSEL5mY3z/TfAyjqZJMV5P8Lt
IKgZaH94q4xyeYfAusrQr+2JxWWX4Cy8pTto3knmvFpRTDakdsz06XaY5t9LPM10g11O4ZzRlKUm
XZGfDigKMNsQJVKWEBjdHJOqJowgooOKhTiDJO9fKeKwBXjP1FHdDbmVllOx4zVxj9218y4EIAMr
5Wg5XyCkZVoTSp5/mnZk1HHomx8IP4uZiiEVPXQZI7NxrYhSdNv7jYZKgiPKU7OmbVK8nlAIrjo1
eobBENcmDUQlJUehVh8FwO1YweLyfjX2FA+GKsqxatxEhHitr+Z3Syo2wBu2gtYIWSeSFio5x+9y
eribzA2KFOn3T7WUfF9YY/Hc08YdWGSnr7jA0Ftp80Av6894hhxad1e6gO5/x7IVsI6gisb7HAUE
cTc2wC9GzNL26LWLzhBUukGKrNh1d0mxmwKnTR5Z3YQKGXWIMjJFOWpn1fXO0R/XPYWaeSbQArHO
kP05sSfQL2DA9Dqwgw/kmgwOzUx29JUrK5eWYs3p98oE2W6q/J/a0UEvbdKYOxfih6NLMtaBSiPZ
nJ+fdQ4kp7iZWNPsMd7BLbavetBq9xLpSIq3LX4dt7Zdd7d560tlLZNvXKw6lX0Zq8US0cYJVTRL
MpN9ikB93jWCgBAS0rPJB7QuuWkg2B3/wnjwcDR0vSfOnYUkjRivH6GyRcliJTK6p7TAgTC2bL4V
h/pbQt60VrwLdEFRHJC5OWif7ZT4lrY1+DuJdHXEkfjz0SwqnfxQNff0zbIFw3XYa/MCrWO+Zb8h
1LWl4ojS1bQ41+6VFLLOM+QiW1lo9FMJ5NOJ2Nl7kKhRpYEiJ4JgN4qoMiAjLEKpeYXfe8YqJhQT
A3JGrw5dMR55kFlJgbeNZj9LEgJwAsWnrpizZp0IWfDlvvw5Szl9QgsAVGy/+OHGIYyn7JwNKW5L
OH7nzB2bAL638R5E37epfLDKrjrNTyV1w7kyDH2aZSC4yZlMF/PJO/aB2N3UVCLX2RatFevO0nNJ
2g/4gMcwVyDjS9KY7pRL97BWf563fp7io+QGdcDxyaXgEu0bEC9dAjm8S30iZLmkmgyIq0Alt1CM
L7Qjq914N/Inz/oS4RM8jqZA1nzhktUZfEpDjtgxYa8IPOjT5/3yh2kIqC/vgL3qs8xjmd2jzos2
1NlL03KTDm5YCt8aWVBd9sk9GicjJBupCjWjBaNYlHZHuSperojB4D8Ug1XwPFE03FqL5l7pgFkw
Ld98znIqBqZNpi80g7BltF+JXckJDZy3sSXgkHbtSf/bN3PYUGLWa4XLY2K3uti1cVwcp5UL+F1M
qLRpGpSfZ8moiF96+KgV/liHraPr9qFhoV5WqxkdWL/ujk6h8zAT4ZH3rgxq499SN7og104zJ5++
d3Q6HijmorYzU800OeLlEgbE5/EZxtaxFk0eWEFzaNIrdbMfPyEQp097dUWruOmO6wi4zWh9tyls
HBMK06RoORy5tjjXd4Igfrnq//Ko4+3/bmbSuNgHhoDPnQXB76WPDhNaQzvBNvaWjXsTqPCWu4ou
A2d4XuUCPM8Hf7JrM52FYKiLXD3LWWYgZVWYWkhikcF4fPPKE3TlxSwnFQ36LQtmv6xkC8FfCd76
YJfSFY0lUiZHLc+xuRegYmEAb0zj+oaun0m1z5ZUgKHQC0sM6+FDQzoai0bkN6mtAdIp9EvJTPSH
kSwZGcWUQoSC4/4RqO+68Afd+Wu2y775ocLlxxIgVoI/LkZTxXtbVlLCZqUmEn6PeVu0g/Bp+CtQ
uFv5eAMALiBUhmT+JQCP9r7cHHTL+7es/bRFRBEv4U+vZQFWd7ZxFVUk4iDKUmXyOFEbfaHc0ZW5
alogs6dUvk8cC7TZlmjYZAdcTg+fne5HwCUG/c8yvGrXlcE+uT1zbRmUmqUSy2Wr3awK81pDHUqJ
+cNlhisf+ulzK+ckpIIGiVyPRDJNU+onysufiyK5i0z8iw2IJ38vH8B2izhRBYTAKkBwBQOHIrmy
05/VeMlDtuDLpaWxJMcHjqjMKPIcArzTnwCU0aS2y/MYsJmBuBxnx4ud6xLTydg2STcWgTakgDPx
Y/TJNRTPmjcpEEXSs7qEu5aZptKADwrqch9wmrXA1jLju8Ty7JsWvGuNNOByfBNWYo0+0SXoldQE
cSv2MnV41hwmLMEeb3dOa16b9P1AWIAWR3+JwZtS3b1YYVSsQUG0MN0TZr8cbRoHBvUh4HS4dFYr
xqLOc8qXEpjvvGJyWOKjoRZMz7L4DhfHlm05cWnAKxyRVBAyZJqxEDUgiB/qKWktzkSuLfxA0RQl
v2VZMmxyWDIrPjTtvg/xRoOyttxtrH8ZF3oVLDKNQvSmH6vMWgekMJumbEFh63gzsvcFGjdtW3oT
RSWhgpJPprCJPiU8yvEw+fRCcg1ABkBZkeu8UUpvCL9RkPWxCBflXtFKa74HUAj/kXBDLsrYKuPk
/W3tCdcOA/jPWa3TFOZoarfTvIkdfQKZCDoTThICTo7WPOhBQjWDgv9P9Ya5m7g7WHf0RXdKOes4
xlQUbaDHfcjBG4qOe5OowHR0MYvumOfJAhih+XA9KLXatpvsjg5bIrR/iS0K3WHRau1QuATplxac
S+3+vqBTer7MJGUDfq0gcZdz+Qp5F/P5s3ak0GtAwm/Gs/mzl/47haZ7iZWNnVoXgFtUnkf29YKf
lhzS194WWRGeaxzIRAGPLS7dC7F1r/uYycY04MaM+rkb+q6brbPpXjDCoE1fujCcCF/Oc6UNPgYQ
5Qi0qKGJLPZd1AEVE0DkQWKoOOu5gXb/A0d7u0ijNOJPpXFe6v9qF3PQaGDVJ8M681cMO0vhHoAa
byzQpDO1eUeYSe65unfGbY7/2tBvPnUquMDW4k7zObpgD3fqE3pS7gA5FgflIgIA8J3RsAArK9Rh
729b8ghO0U2hPQg4Zog8BZSAho/HhSJaBi+9YkCdL+I0wK0NE3B/E85ELlVKKeVZfcOQjKr/rUKO
60dund4SQPd2QPythcKwPL9THvJH8s80EBb6xhZtXlZBfwK9tok6ybyxyqSwY88/6tOVtn81EeBD
DkVFH3Lq6oKMblU9MnG7VhiVr+WyYNGyYKPpSVvFnyBQ6aLJqp4dzGmSyuc4n7TZDT2v9b6J4rbZ
NzsaLKOdf73qMtvkNX8tY5yEko6KWCxPokSUs6xcoIlzmjNXuTYWKdeV0BnHENBNE1Ml+6iRfn8f
MaArh3vJGaHZH2zyr+v2mYaeCohtL0tJzz1gPIZBxxNrM0kFQUtRBeDdahSwNXwRt6W21zr57lhu
dKJ7zJhqzGpziaWKd/OQLrtysFJmv+DQ3dDY9kIjJOJtgqb+RoQYYbR7C71LYWLMUDRDKFkmJJ5r
edqFYJSzWAAGNSrfPc+DyRSZ4dSunRzI2nlXx5Z9jdJQmUdjwrhbJHfIFOgN7hPbx53nLkxhgflD
3itoRkUhqhsH69uzzlN0WYOU8mANzMS1GVsoIrHUfx8pHAgzh6UmNeTjYEkPTW07Yf7i3VLw99zn
Jw==
`pragma protect end_protected
