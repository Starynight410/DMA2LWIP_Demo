`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Jo0GTP48lurGV9QI1c62RTUP1YVEamMz1VZFzIOsgfj+B/Me/Uz/+TNhvOgX00Boh3rVDWY3miWC
6dvD9WUK3Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LQaetkHlTEQ/O2QuW4ImDf/K0WBzrX60Y2eOh0Fzlit7V6+gYpu/pdjpcV2iUJ0OSkPSJI+Mhtnw
My00nmvcw7hr27JQMftgpSq2KJTPiuvMTKQgaTjH7G11dDQzZg5OIfVuhiEdrvLjBL6ODFpLjnot
+wtza061w0h0SULGF8g=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e7yz9u7SkKHpUf45ToebPKpSB+7SYjKyIPDWMVo4RpE1fApRY5i+m6AdkyczFN3egPL9yuxMUBQi
B3fcWe1KL481lABpqgSqODHUHO2V3VOpcYtVbs+ITdbbKzYLqgggxX2OFaFxfaKpm8KQDKkYwb5s
hDH0bmxkegiSbK8/6cCO7THsM2QEi5MCtiINLnSFKZxzW2n5D4XuM/reG5kcwrmcvNmgwL09iDms
zsLNFk+KlTwGLQ+sjNp4XMp3wRVy8au+yG/ZaAjv1SaonTr0s0Ktoq7kpKzzK8Vdx3gxl98oC7lG
qI6lKENHTJsj2Et1sJqARwUVTfXhIwUnx7z+eQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YUgiCLqe/j/NhPlORdPixdVwbLBtEL3BY6gCgf7tGi15P5FTCSoEIKV1fMOt5n55kUiULz6ixyOx
w6KSNkCTxNK1tRyjWlYPNwh+30X1DX2lqxQedujI8dEfW4TThaFzjbr5VzZ5Xx3QklpDtemVWlfc
v+85sRR7dpK2+yz7JHTpwsBUmUIz/yQuKTPH3TXkcTEtK3SDtuMd9W57I7EJRQs/QWb0HRC1gqri
b73Bznz/ITOHvk6hyVhz2IcLVxpPIWw2SPni76CtRBGxpvEkYBsB4Tb29iojsozDmdeCBCdMwy/R
z6g42MtTw4HdwvXecIHU1Ps+g//YLogOmAG9jA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
m7rYtXUavsevrUPbAA9ErlXCOGGk4fAoeRrucNOvvuTkTuigciZtMDGFuNCCP84AUenq7yf+knfr
YxGJdpaWbSksXpHqc2OaU9JxiGbOYXsVLB6aaIcsBViJ1Iu9Y3dsxqVRuEf/+KOaUoj9MgYpzlBd
dGJCSN02BKWDuiELCvkTzxH0HkaQw6L4Fs4eaqtvZO6JC37ps+GYsLvCsUVOUrxP3ZXffR/5rO+/
r+Y7T74S//4yP9CGXNTnVBNea7FKmyEzggzbDLVXfwg7DC9jqBdVLhJdArtJhH0AWfbyCLDAfF69
TIFn/nOkcwqHGmFmfhdLuMOHq1GabkUC03gqCw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WkzTVLle3kbJDg7jpvQ16rMwFjgKsN6s5VraGMgY5PuWLmuM4CseW8hGJcsf4WjZloefR1XKRkv+
EV0MnXlsj7dM99Z1mYpSYEt+FSSlVw8ZrTFDfAXM2tVaQ6tHWq2thbcjDszMiCZNwxeaVwffojNF
dPRWtPW7gJ6hRMZJ1oE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nB0LvvHetoBgxBsMSEPN44HAKokSVtsq+whVeE4wsASFbqJ8K82xM3hbmxu6ZDYkwRj1/AOA3HVk
G4ilfKGLy/G7TDbQDfRO+5Y01cbhrcP/GMxbBzv8olyMaD/JTd0uTncjO8AIV8tUE18Kj9ZhfRCb
zatytXSeRs9JZ1gbnMMyuS9DWHly6IquSzk4ICOoWWjyjXwHRFPGPkYHKeAKIXuBgNn5YIUb73Bg
ZfSxBEDnDG4lR9r5BsXVWXPmkRPzzmalgCEOM4dNamRFXJG6Z063apEzsaFADjlPswBxcO39daPt
PO0nWMUFnDtLtq5NhL5JcY8vaGgEnfVUj0929g==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kx2/4FUG+WgpOeMb3Rbb/cih1lc163wBQ4vKkckklmR615Brrk0uvh47GWx5YPIQIJ1dUYGfGof0
suWssmlsLprBF4iyZ0oJN+doxvhmSoNuyqNtF4sOBh2mA2fEVAiuuRzdRQMw/lsxuNxU5tTeu4Hq
m6fseqlUS4i/DqAjB6NT+vlMZPYsrIaV5xH4A+ZthsSp/Yv1VhT2z1Yf0I1zXIDSJLePBat4WiXu
ztJa66W8SRYkuIFjEUecZElA0JE2MfS3tIGvepvw+Jw2NqcpRNOyHazWtDF1qGPoplQ2+iAwhvFE
swC4IvCafgzOO12FbZwI5Wi1IC0+7hrnR+7e/A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
8GvLC41uBcFwr5Ki5OvQAwh2MwnGKfuE0FkJhaohC6KDT4SH9pKcwnvFqbHTm7H+kxpfjlg3NYlo
R8dPW4XArskiR6Di2uUoB/KHQZgA9Q3NGeadX6Ud+7YeOvmXZHS9qWcWSKB7Tg9k4KbRA7CJztYE
5fSwBn6n2UJIVYg4b5prEiLhaF7+80O6Aj9awHpU3/4oTqslJrrOc8Dsd2Y12sXITAkhxRzu/DxG
fmOGYrh7sMC7XdsF5nOdO2hyWDVnNQJgv4msDpn/EoABTfLqEdtbM1wPYA+bOE5VO/ox9n1YOjFk
6mPRudLGkx06I3ng43nr/g0r5vdEHZOH2LOzmTRLDM35vOfVLM2krQGukkS7/492CRrx+Y4QHVl/
GBroOBxcUC7n/arBAspG5NvcKuGifZw+yQpZK0SzECoTuxsXXvsoiwc8j6SRIhaAgTqN5ZBEWxi8
FNVnK5S1778n5yzbh25Yo+ngzmO4c0rx5cOkDGRBGD0P0fo/QDXc2iB9IeNitVd4t1T0ygUvERPu
U0K4ezCUuRdDq2P00mJOO9dVy7tsrttn9SkE71QR3RoNDh1aba1FUHDhACDebSBl65J738WnOP9N
ddE2niqIm+h2ps/CzF4XFrGvyYEvpr1gzwiZP+jlZVCKmDExxS2/UzhLqH6wUHYqW4ReGzrCpQ/F
7BgxbHghaXUgoeJbXlUJqwzWvsyc2EhKjmCOLeEplP2J3HFjJ0byuR5XNd5RBprwB1eLUNu1n9oG
o1tBhH03ovU4rQArf/n8zyeJLq9i9jsyVDn1NfGM60iAq2k7aG5U47Fqyve/BKr4UnVBzDY1YT+r
wFoXYt3oIaclzYB04Ku7l9dhOxCk5fdXtxUz3pVc4cTGi8pgu0vODpTwINXMrh69MC6ccZe5qseU
C65xRXP2Y3box/ZVst2BHCj6ndKCeA7CSe3Fj4q+uFuCir91D9HKoPUXXn0WmsZOFQ8ad94wEChJ
6i3pQBnIgATLVYWXeaIhScprcvBsYmNaRm1zcf7A77J3pAAs9+xcc9Vdl8iWhVxGRtx5ozMV0akh
ILjvvOF7fjaYO1eKeMvVKnjvaM7ExUKb+4jTKBHvTSCMnNn+5IRsgGaVnApRW23JrXJ7NzggAuBN
fBNpD/+ek6BWsuK17K7VH98UwG+Xs9su7zjYKR2QaxHMtqm3P/CLXoN9An7QejmJfVrVgx815ww8
vKSg4T/idC5X8Lm66bYy22PAEWi12HUuzp0mtTrPlD4tUI+Wj1bErfcTItJyzjVAf4QjvPoJ7qIF
+zN+iYlyzv5thQdPNUtv/3AykJBs/UWb5+dav02Ry7ph207POxYSucq4m9m9KdrkCMJE3E8Zqkhl
A8L+9oq+wf+7BaL8Iss2U06HZiXObm7r785Pg3fV4crnUorleZZXDQ1jddLCZH1neDmrNoPI1zva
y+q1OAxO0IgWNIDMJ8rcJ+S3MmS1w51o4P+Ja70uqIgmZbc3mA0+IQfUHR7hyQ82K03CtMRVBLdC
KeJ1gBgTyYi7mPQ2Pl1/LSkR00DC4xYE/ZXqe1Rweite0CI2DMdu9qfRCcoOplzLfPMATHM7EiD1
xVYObMfYjxb3adY88GnOyCarV76rF7D+kzXBFdhtokAPgvYi+QQiijlvDC9LccyLoGab/G9APOye
PENDGwlQ/4+v7EVRq9YOeu04KJPXFA8o/HZjwIi1nrfR3PagnaqIVV9lv3NsIraV4x5Jz/OKM3o9
0mtaT7GIrALTbI/EbPbxF/DfbM/1p/S0XIc86dO1DKrPnGfvjO6tf/eTIY/F/S1rVZaLoKCa27sO
RJWmP9P7aOA1qtAu+Pe7rZJBWBsaG/PEh4T75JWUCf+9aS5rHU5WjVvQt4JvKRNe5RAGSQvnG7oa
gDBesjqosrdjDW3lt93jrRwSKETKwFxGyfDsm/jm07WuOXZN5lCRdtMVTKgEINV5qyK2pI5aSqGY
qpmoW8OffgJ1IPAc/MvgAxKLKjkSz3v4fax9R3s7oT8rMqkhme7km8zYuo1NGYzHrxxDfX6Wi9H+
vfspB/fxBWzQVq7iOnk1/QYvIZ0Qel707dWIAmHDhG5q+acR54E8bBmfTTcEzDdAeTy/88FWT7zK
Vec8QQADu7D3cTgqA4WDPQwN2bMQn1ghvJW33pSRGXo8SwkW01AGPCrvYpygag03YgWoSbVSgipu
jEUP98pm6pvqEwluwelU1YusV6v2GyLgtXryR80EcqBFx2mYJz2/Ib0a5+5f+PHq/WoxJPAEkBki
ZstzXZDYw+Mv3IDIbJOEhU5toCFs0+SRU09Nc2G/q9AL4VhLkEg/hOUzueF67TA7oHvJMCv7n4g0
FKSpHA6lJq0D/1ecn9wbgbAB2Ip14obKjQCvOjaxpqMr7MV1tKlg+dYDcOkRFYIxbw7DRrR8Rpih
mB+PEvWixj9Ss6xG27u9emO9mGNIieDaGxbbSYUKcJwQ21gS6upjlTieYQZjWsSKuBe0PGEPWaRT
6t2LOqLm9poqYx2lrU1IZvwK715bcy8MOvn0aRedwfAa4JkQPYsFkIeW4p8pv8/67tulJD5klFJq
CVxFpHDNV5cXgAqCBT2J3zy6gs0kpGCZLqhbtVGlH8ZUmHE7lNwlbHfmyrvOlUaOETqD5V/lZ+Yz
w1kaCVOgD10EyprPvNiZ7/1ef5w1U3NMsZ89wwmKRdvFst/YIu5U17MHHKzE144xD7UkfYpg5sA5
KlvHSGC3X+g56G7iDStJerS9acu1hHSBbJeuAve/KEx8i0/hNJ9N4BZM2gz9agoVsTtygXCUSMON
prLbs9b/w+EG3N+fD8i2d0aE+FZe9QCv7IPfReSy5ikm8DGyj0N+A4jbaNZodk3bimCKtMWkta9d
82/wtyMLpi4/rHWuDu3lCzdvAIXnwoBp5vA4cSoh9DXrQaSf5lQfA5UirmAPGlESii04qSIVegcE
FwevSU1w9xI1sKrf2LPdp1p+MB72eXbTQY/5WAmEvohk5O1tppJj3+6USKsr5Jp4sh/zZLVb0b/T
tXqHWrXCrtapglLR1cUx93ixrQqg5yRd9olZiowOd+6CoMGFZKjW5Ny4EbPf/LQaWwYYHnyK5+87
4oU1E8Cx5wIb/5ofVXox5ehqj2GkrSoXSdZMAfGjy9+/ln2pzKWT2FwqUJLjOP+oqsRfKL7C2Qc/
9Hxh5hUvvvcjeSaA83mKfVzB6gc1pR3YgF0QyHtTkn4tEJNajDGxmvwY1QxKWXbBSdD4mahG+nhL
Jc156bDFGuH7y/gpJK7IKs3IdQHiehCC2F2q99IyclmwbUkjiR1TaeRFJk6IjATpbYSxQOrv0YmG
WHanU/yfgtmKVcqDq7iPakniPxBig+Ewo7oNEPW5iCkcJ2j5q9i+m5ljiwAqJEI7O/WafDDJZcPY
eNbLEOIhOhTk+WnQwE0FoXZUsdjqkoGuC5ac2G5Rnzf73lNF8opqwlkj4CN3rkbCHrTpx3wBpaQM
5RMbgloaGC4GUK++FQdmvvYmNHSUp0mmQIW6EZz89NiIdNln100hYpG9SqTBuErAeqORnF4/V6Qz
akNZvLKFM67GQZUjA83SgBQLrQb+cFpcQtjHIFAFPabEo7vfHE/fV+hfG1F8xs0fP69NxBG1F67H
N3WAYiXKBJXtLN6Q5lG44OlaQ+8H+CujFaQo69elxP5/R+dN4fdGlLVn/NKC8ZqmNin+QWa3+nn4
zoMH5kLiCqE6N8MhZpdqWyIwkJrF9kA79h9iTLrZHGJLTRPKuq6KaiNP7ZiFX1L/L0fwoc8NNMfx
hcLSn5Dj2mmN+lbMng3fiQ/mSdju1AWsYkt73EGdWRSyTtbYffB2J4Lk4jzlCWggj/Qbok/fy+iq
wymDHXB/oLOaV0E/yspa0vqGkD/LhDSTSHniOn0gALtOXGeqOwjtw+7eBw0DLzC6Jmn9d65IQIg2
adUOqL/KC/AiS/H3bkuZg9WbCQMbjPKGsivLTEQueeNm+RNrY2cnIoDlwQbuy+/PNcrXkfVWCS0I
KSNctBUYFZnsBs+sClYJM9VEgZVcGVvHs0LMDzI9kxXtuTXhIEWypSd3vV3zJHvMzKGtipAxD0at
dvyg82Ls2w0N84v/m/Nc8Ar/I3Y7AMnNySgt+nD0xAXStvHcznxdMsXwZh73V1R2/K+WiEsxxBCZ
ekM1r+DI22/pGQqHyGBq57x20yQdGxDK+4r0MYkQFc34QWTEbBxg/RvYDtRQJY+ZBZfkd9VnDMDP
cdcQKt5CqKqRMGGaGHpnUrgBgwx7OutTDDrgxXC+tk3YaTAlpSqFuxqiSzEshqkIOidoaYH1xhGe
F1Tbkz8z0Nbrd9IR2Yc9AoT87W9BFL4IB0OhVSvlhNThNQn1XplOxJIdDstCisHnlFN70b0c8ivO
sFYpcybUWf6nDDxT/TDYpzuK2ggmeXboCppeYpepxKs3+Hhgg0kr6dQbQxZC1GN2vatmIrKZGFk8
5iuhz9RGDzx8PpfUDY9PLWhDfi7bg3UM6QW7Ho2kseokGOoD63BrBb6dBZE5Fd5+JdmJ5vmo5Pv9
f0x5QUKzds/i2gZi0koyb1jsd2/XfbrEJO6b7UUVhRxY1X/D0Dqqsa04TpI5d4dma3ojzbphoG5u
2+Ayte8cWpdtXhgc1p7g2/ABQJGQm18//1BPZbMZoah2Gk8DnTGhn4eptbZPHG0iMr79VvhnI9jz
k61ppud9EvvvqaHJofJOkQ5g3wDArCGzwcJRl04NK29prLP3xN1TJsAon+X+3S/GUZaZK6TC7Hwu
Hc1igrZrGrw1X4Gkt3aHr61Rt4PjEbU9hFOyFZ93VnuF3N8VCjLDP69yIatmlQPuoD0+NGfuLpFW
9sp50Aq0mqNd6i+fXQe/kzEktOtLYibYWt7ISC0C756iOFuEDTV+FYWjjjB4NQ+6sykfk0ny4nEv
Eg/k7PXPof1255AQMosG+U2mCALptwdLls7smD7siNug9+IXcxIzUcGSomcCPvXDoWh9OJo+GtYF
BN+1QIoFeH2rama2+ySDtqWmARcbJ1yIEtxEf/sjUpCvm5/oirGqGFDc7Q2dcyaru6NJvzcJcdUI
Yz9RIRFoHshwD2oQO9I0+uC0129I665piaBbsdNTZKqwF3/pvqGH+1ink2b+4Ydqxx+OoNRrc05F
zvFU7W4fUVItuGCU/qN9GFnDvuUIjJiVu014DO7g9gp23FfGJNyRzvRz6yLHYYtgVrjBrh9UltJz
/mu8R5UigMpDhI5fEg0B+yfp4/qAtyPKMROh93xyJ6yXDvv2T5K8CXhqa7X5yyPOchq9EekimJKL
IDTKQewhGIOpCWOLQnyFN62VUltPPlkNoAs0rLlrDDGeMnRRFwbvv/gQ0NbOKqwuoUrQ65Pl+XlR
rspgGKMmh9TBm17998dtHKKt0YUCxcdwjqH4lurNQqu9T9aWyybvF9G0Hh642JBamW4JI2t2uNob
RaC+2Btkv7I642GgaDOoM/KRe7XAaACZ2qNiJk80+I6wLa/GtWLAOlvEgTR4tl2776vskbdynD3T
sw636Q9kQWMocOwPXEgna6e1X8B9pCz2FUFwhoTt6bufgK8TltHbYQShONoRFO3J58+hcrb5zdwX
BWCIbAuJ4ChUlZ4j2edw/tpWV/YP2291gSFr1FeK8Nc2jeo/C+axf7UiJYsHBJuithLMG2+XawO6
j49mX5G+57+SFxXqj8VKiYF1sTBN/YBlmDaCkG+8j5t6lRrOLOsc4FMBWBLYbb+RbIxAaXJHlhrx
v6K7KlCo583lshVLgn8EKXxSwKuU4nqFDqgbcPNKadAkDAlZfJdhV3TaXCn5N2lEjRp2K87/GfuN
xN0fU/U2SBCmSeEkqABCRAeI5Kfnp8YaqB5TeBVuXzKG8dnJdeIR7+WveNCsU/7t5eil32nuFzu4
jmmqk6NhTNpMv19LDB/S8YOAvMik927NWoIqPoEEeEZLbP2fCes3P3iLEgXRYMWWxoxXqthWLrgv
uzSjvXBOACf9TdW9ps49KSBeXEKPf+x4iIxyPAz6bVPxJn7QfsXo9urCoMSeg2d/ng9aad1Xom9B
R15fOBVPtYp7/5xohHXgpVABWWvuuhMw7NrPk7OKzhMce2nEix2ydzZYgo51rQyei52kLHkAOjPm
jpund3BRsBpLjuLlve8BHu/M6UYHDKY/JLLBjr4jmQ07AcKLThdGZTmkLBG9BCsg5yskniR9q1QK
S3HJyIZgZ+hca5CMGevXME/AIC1NU55kgiG5tpjFkkZDjWCV2Bl/xOuRurj+Cm5lchk2PhI5dRNM
Mb0r5+03ttc975/Dd+b8KGzHyVHNHrCz1+1DSCROvO7ddFUc6tHmurBCutkiEoUVXXkWkkGCETUG
eHOB5RfNhYCuxIbLnAtHU4Oq4JGO2WhZTAPppf96emv4TD9FfKgKiYKUDnjwE7DnvSyc+uPGi0d0
rc+b2/ojGXS+qa0777lC4h27j0h3e1Q7FhTu2s15o6saUpL0mEuZS1z+kUX+bP4r5lwiZ6Ko0LsA
xyfNx2SlysnMjODBrkefpjCXyJOna5th4vjcdyV75N/KgilsXIreq0AqL/bXJuDzHO0y7Io4V1xh
nzLeSEfVasj0mq3uZHmSVWTbIPCX4VGQOV7flOytst2h5Nj4Znpe7qaQQwjHk22a4u6uPledgYl+
8ubS70bHZ2PrVdyS/SJrbZPtUINkGDkWbQbaj3qXVQ/A8XMNhpeQNJGz/FnAGSQXEWqn2uZWfSZ2
GHLwoq3Ns/TgkkyCor2qAXzfCK848vNEYHj+yHDcayTc5bMxfDplLfQho2OG6sT8MYF6g+Jc3C4v
FVrzXyQ576ff7fH2ksTecGJhnRUGBFXH4p9h2AEQhJ9TbJLdUfYdtXmbKC2scVMEVvGOTuBKUb67
SWdyK4WgI1bAcdGq8j8ct/IFMkvNpp1iFEQXyru++PD3oSAw9LmLWGL0XggbxdQ4BXAV8sp3lOuU
Pv06CuiCBwh2E6opMxJwcioFi+MZA3t4PZZOkNKFrFPOO/z97sB+7HeuN+z2aWZj+n/KloX17X23
//0+52MCoLh3MIQ5w30CpVCdAUmY79mfIA0Nf+fmEtnERyIg/ye8aMujWfkuzgdq0ZvH6gtCX6Vv
Z58v7Bpa51I3AhH264GiyfTm82F/7jn53WdQm+EP7QPjcNZS2uV7abOn6OQwerXHduEQeUJFC5d6
ruDxoUG8NPOoLxV6h8/q5U10Z7QyMbcQGOSi9vpCfY/CiD4nMyEi0eufWnMpVpqdrj59RbuFcnhA
rZgNPt3MSmIRKlxmWuJUZjzKUFH628hchetLR2gWvWnGDFW9ZlYctLDHbA9WEOwjhKFEkDcV71Rq
PyFscctwrScGWhCEeSS7DLshMEz5mcO41hLnKV/f+JkIS91zgFlabHQkuiBz+pMGur5vRHpkujRd
Z0eRVVhvVo++XW/0pj7Ct5q1+zw/TyQWTso5cR4MRgNSexTsXg37C0ViUA2IMiccOk0ZVwfPI0zW
Ggac4ioEertckpMAUmLKhppYgfOYWalJoWdBxIUM8+AKWD8KSKuqZ7uIeC7Bsf9q4s9zKHNKvcWY
Xn0uah7MRI/a2BUS00S0X9MAqGszQ8aXo9zOnsqCqWcBltPxPZ3AMZwb6UH0xFQPKc0Znlvba5Oz
66Y/9dvb4ejNKpeA4XKGomZzK4xdgUZy7gvV1ATeA/Wg1bxsnJmgO1uj7LNT/mQ8jbc9LK70ArNc
IJlSVt0f/YIBv3XpdWlNZHsN3OpU4aaZff/BqsPq04v9obb5Xi6lMEtlmJs57nGFFKXeu6RetmeE
yxcqlA5JMSEswR3LkWKChl5tRHYybqM0ZKFgR5UiYXQ8MoIsJjRcUeJQSzbKIiaEzT4fbdjyI76M
sVQILG4SGYxyD6Q6qcbT25jc3/OW0fUpkNU1XX2EJw0LoG/7FzqX2FAmmK1XRlQxglrOTlUyq20M
DTDP6zCnLqxnqV+d+iPnOgkvE7HBIOliX3YjsOLl/bkzurF+vZKCqWGg2ZtTUk+7tOE/ckD/llOC
5R6gmCubyBB2WzUAbYfGqp6A2+MoPkasrBlgVp6TrhqFI6hxmxGRUsc2wsu8iZjDo2Z7HcjL0KxZ
kGR1Oo9i/74DI+eequO99CavT7AHtW/XGtSoVZ7HDZP6CPOkmARKjusqVko9vxi89LLfV98YFKYX
VCDuAvIr9EoqYz2YFLS7hEL7EdOiImJumFwoJNPO9JKX123f9a6PVWZG32rJuWssM9wySspTUZef
Ti25Li0dBVJqr0yXCKaxEe0KcAus4PhLC2+bG9kkF6gtjEI5tK14peywAw1NA30ypuDoY73GIJjo
krwB1+Jn+ZLD+VRWv0wnvsvkNam2fnVuLD6qy456u/UgtrWgSpYRqobFeIDwQpBIp7KIYcSYV6Iq
Ic/ZkDV1FDWXC9lSvEPP7IyAtrEVZ7Q6knIZzXDTFmRdE1HTH7vO4+wclXUId72sJvC4Vrj4qKdW
R4WMYXOKxyFbG3CtWubaP0BtMC9zucypob+UhyeesufJVI0v/L2A5kyKdv6/Jz6m4cfbtWp6CUb4
ADi2DJ0oUdBWjQ6kExudDgG0lJn56IfBCTLxXxyObW479v3gj4ZP63ffNPx22mA1qs/l5GLfGwkb
8PyZv0HFzUIgmsfGeVJjwx/PKdm4slBmuc8l0OOKHSaia6QigbAOqHQYOiarAaWXaVUjIkM/LrgY
lnGJBCZ2zEGsXuydqFCjlENtySRiCW37+cAUx1KGQZ2AguDFTWrg6lr/thRmqSbWUa1UFzqKM/Tx
i7nQ7Cdcl18vqVGLYlIs+nGoRc0h/NRLJBcG8NDfiuuMZqX9WroFZZSHAPhenh+dCtM6r5kx8eXr
9mO0Zvw7Bd0k8WqnfaA3AZM8+MYlUAZJUTKaug9TPJ7YOo99V4ce3h3TcaSrN+OIIrp5Em2TDKzR
CJb9wncmIhHksYA5TqjMOwUd9SQOwzHFXd8QGtvRB4cK77/kds7JgjZhY8kspEgUXOKX/2Jz1eTS
sOycAkGhMekZbFX9DdERC3SnRh7Ipww/K+S1veEPKC1Sip057UYO+6jHeUj1FtWA9OaGyFU98JSQ
5/Uec02XiaKbCDdthSHvsP1ebwFI4pC6PjYQZt/K9HQcQ1rlufj5NNYxT+azN9X7WdDumiGKSb0G
jEs92fV+WZg/gjIc3ZcXlJda+s8JTgj/Bt7nzs2UnDeIoQRrSRQdDThXQ6x5GwJyZbLv1N5oZN2F
Y2wrS/1y5/z2XkSpgSOA+6Qj9tkiCXqN4jbG3CL9UZ+pegm4vJAJzK88ljQK5swkXt/AvG/pA7wI
9s7FN8bcjNqDyL0lJeymqdSKbv0tJTtnFgAjMUfQmP8Y0X7H1h4l9WRAHUyJWSNd4brF3QsmopdF
lFPI2Zj3BkcNbFCxIOD1Em3zibEAt0o1Nd4kacxiBxcj76lnGPoESM9VGktRkGOezOdwHadrwPkP
svIFWgtWrsdTPKE9ZFX57b+lcgTZqE0BxU0s6zzvuDpJGHt+HClnmF2z85zEkRcHrmVqKWuUUe3Q
GBmAHH3UrWmjxdXOCy3TF5tidLHK1Ip7ve7wJRxOWLVLn3vc198BPBqGRSDlSEYlCTK1DLgA1+G3
B+zalVKPhzVwFD8YqLwNTXLEoCssPHWmGK1FdRH6RRwKFSp89UE6942N0odkBaiR1alhfibGlnPX
jRs4yIud11f4bBRA6EJLLjS9Xm9PDruNhvgs7Cv7PjAbUwrXAaFSRJ4OC16jbtPAH/YxG/z+g1Gv
JxrgsmV9XBeBsqxzaSqOovKSy2qVSMD3M9+ubFzA2Aj1GNcwMhNo0KvjVqyOOYoapUvd9L9hx7VQ
SU2agU5b/M+WvmGW3jiLgzpt29e5eN3bTlifldHCrOGHDRgBsoGDbY/ddHVV7znhUIe06wS0Z7ei
mQwob7GVP0Ke9DVNXBlwyhl+du2ohWRB0OydS/eoq4HRWGu2l/0todkpLx0jcEnKzjgNEvdHjIll
+DZiZuq1jR6dfZZQ/furSVloeL5nF0F9Kps62+9ZYVrdoFnB0/Mrwm+MfzBhPpPynUAw877f4rmg
rjAljLKS5nWBUi3u5j7eW6lU86R7q9ZAmCY1UpVGGn3w/gO4+aRJYpgkSKI+am87xEs79PZ7B25G
R30pqgvvVcAd4ghG5n7lL6c3zfeEWCOpYT4QKR0pTPflPZmaQ7R4wznqsrKPeKyVFTA3CRawnNKp
qeXoEHmdEwQCCEB4ANYWepK50lCDD3u8DcOfirloMjv7jc6u0l7iCpAgNwnP99LKiizaAeFntxeo
p42ju+yGGHLxwdkoy39IHAOYtx2urOPTLW4eGUXSabVWb7yruKau+rVrWrkgqkHD3UvYsa4HquU/
w3iaPBG85sl/aRySdgeZvRt12ovE1V7b2wdpRS/aNRjsDGirUrhfg1kCC9zi76EXdcNFpuTAQ1BF
xw88Ho6qM+lb8kQyDmMaLqJTKrsSlhiMKPyh++nWv5q9KXWp5J2vcL4hKFwAeyx9la0UHv6jY/1r
tg/nuzBGAcMLh7fo9qm2pqZzI9XIWEYozm9m2BDMaU8tqbbxm+/nrLxNSe8Hj16iD1TGqgWjMqTx
ZmZJTgvw1Lz37BVFFmhyb1dEYjaIjYnPbzqaeOuUnMRYAqhrmw6kF+KxxLRK8GPRLCbdk1tX4B/v
tvrY04EBrkus6uxZcjgO0H6Ii29cJGFJN665/LyAWl38IVxRaEnd1+YcsmfW/egiqW9zPunkETA1
/xG1i8Oh9yWB2QFE6TpxSzPtNu2pIlQ7WRJfkO0ja36zKmrpD9A7Zua1mJc8x/TTGLjULtFFjZK8
ar+FFA5JRY57Rf7Kfu+cOf0d8y2di+zj3S1xpEcnws2E02CwtJO4G7GkTNL1Nr2awDNpArGOqADM
SGSdWmGya150SIaxafePxz4tUf/dqmhciceAgr4JDyYZhNh9L0RHwZX6Z4ibLpDD+hMrfs5h8Z40
4CVb2HirCPvJKXRP2XyG3VOdKFzr3sUNJnFGXhI1h1LdH9jyM2SvnV+l3feh8XgwKpeEb9ua1Aje
UlJjnc5P2AlMEjYDRsINWwjbAqTaHRmeQvwybeD8Gfj5vsaY5wUHQz4HhWZVdUXRp+qPdiOIpA0t
dEcGqLgRRLqrda55dCkhVL8cQC6JZXAuxb2Hjiul/J0cDaAZMn8Xo42MJICTixG6OBhvxwQHF81d
WO/dHfoAlfaPZu62v9HlEz3/XOiflDwEzbdAjFqIPy9TV3Dh4ZQS/Ky0ZBxDDAYKl9qrk+cPl5HC
LeUCMW9wqAiVgOOQlBbawAzdipu4A48snGI9VAzhZ2c+MRugE+KyRlQw6OfM9XHnINDQsGst2j0l
PxcjHL5cqs47muZbxvTvaSXy2HPSOq+j2MHtdidU828irMWQkp+ZMwOZkGgdZWAMCxOV2DwbcKL4
MKrRJFGtbnrZaFIVx5sxt6QeTMCFsP2e2xgKnVaIfIfYvuX48oXNOSq8Ximr8YctnSw0Hpo6DGB1
NcuDSsV2cQgZ2ZuSOuxND6WHQEXf+y+D2cdL7CPKyHKnOF9yS0iQru6TDXbAi21c6mSEDdcfT4Up
kjZuUli96saSSoE+//92sP0WOnZB5FhvUnI9Pv6V9Up/EbuzLjqM3Dlbq2EE2oyTZ2QKtVQUhSx3
RfLiLSVZAfvWszfvB+UvVVMn1ubuu4QJVEF0U5WxBkYIvNUX6TbbpvIsK685rGDKpNlSoj8W1chQ
HKdWL/IrcSj3hnbNnMkeLUs+gaYO5uQOKQh3i4v49QRfjZuAXUoU1hgQSJsNoHsvL9MyFs7CYFs+
JhpXBdm/SfyOMZf4JwgzvXqVoL+dgwNQOfJWbmF/EbWWo/pVi3OO3jCLh+kWfYWxuxJL0bLjcpDX
a3fY9KWokFMUJAcI0mHyilhcRarmb0zecaFbX7iOZ5obETzjLs3OjwHpfgg7p2K4y2Nh05aWmlr3
79TJ2RKS8Ii8oKe6BhJlVsHC+1XNqJmICHvzy7IKgOMeETkkBf/Vj/7OEVkJOM4Me+jGgUWHScAK
n0C40PTLPzrb5gsvwEtsWtZvumbFOvt0FOlRzlSceGv+mtPkmc3exkeeGdc61j8FAzGpfgOZPpGB
rAh2zwAdFtE0FtnQ5Mn10yuDm3Is5cWnEL7120i8digoLfgsISo1v6nBri9hQZcKU5g3SDdXVnhI
LRCPe9KvKBF7TYZc7VcYHZge3J8i0oCjkdH2tAXgI51U3LTPMm+HumKZpD8uuSGnf56c12fPWL6N
sp3EWs3GE+7w0NUh/M0tSs+wAL8C9A3SC5cQuXFnN5HN2EzHO1Op4oFMGcRak5+m6CQ3K42rEYzw
bd8i2WlCkH2IUfhT+QwJy4ndhoX6Po0ZAL7u7XNCbt9/RtnhQQlB/wlhVWLCSidfhXwATt5CZ6x7
V+mnrZzgUBwX9t/3d5N9Ivy2NYZ6oqHhJSK5kWR5VvbVk4HELKCi4FMB2+7/DothPqX3UTv0i4GP
BoTElu7y5buK+eAsUHWh7Pis3Wd732/TodTmM0gmfl2u33qzarEdjUWTxhRbbbKmHs9b19smPCys
384YM+u3LSRYs2V0FppvaahSXjdqFDOx7CNyOekHbdIxV34ZE+gFqpzuhsg3MOWFc3YKWfx4XfAq
bIlpzzWHhNgBTBy6NsZsuGDf0wA22u/94JbdAymiRqWi/liDI1bfc24QvLTCLcMLKjHuxw84zCTR
65hJJ1ZQWTiPXFt9W3T+Hnggvb37VSG/dRo1N+2RQ5kRAKLg1oJkTEi5rOL/fJmUC/EgrQqjmiWj
+8YTOH6nGk/xoejKrLD6/rnnLJ/qE2NriqGcB/EWnpp8zkZyYZGQq9S81tvDkVUeSPhF5MK4dB5r
7kkmzZIM18ee7nBNAsozn7Dm1Cr6xvkud1R1rqT2Kr5i41Kw6a/cpCp+5NsouXpNBWT8/QNPhnVc
kFunqTddL/POQAd7gPPJFCILHQTPMr0OHqPS4qtOuD3Fgy9s/jOM/7EC1xjUSeQFuFnnknxhjQuH
IJ9Imp0ERX572qF33hwCOZVgGX11Z1AHMAlq6ccNVzEAK2fyTknkdUYBQxsdw8+FpWfo0yGfukxb
nhbH5Dw/q41T/hYpzFfSVwcWtN0mqBxIXSh6VntORzu1iDhYhmoy9/+YIBAePtaEUEMwCU8yEaqT
muTBhMYYo6nZz1x12QbdyDnFLY/1ZkNqthKX6RH8OHPz4NK/pldUQ4JOndKt55JdVH3iJ6dS8A5i
5sks3q7en93QpmQxbrpJomBUz9tvmeJBuDZEdvbH5iUB1O7ZCCsapiXE2MKLdeizwdYj//GtKj49
+P0EQDt7vZAq5GwAzEhJtVlWv/TYyHVGcsvakA4SCh8bdaLuO30WgfLt4ufiIabg27lvknz7w8qb
66XQ9XqHFpoxPlnmkR6NW43kBuspoNcgz+R9O+yRHyJ08nL0b1f8LaJavNpLZPJWwYQywQAAdGhw
w+lz01QCZdkYKTVGeMzD5KotKMuZfstasz53ZSgbCPbKpnNSLFZr2ydiPSfOaUUizUXLvsDyQ+Dv
HxGc0WlttAnZERLJLtwqXyFRZhEpFotEn+SlTxgWicaOee7hFG9pYy25lwULitghgkbFOTlR5MRO
4WZCenEh7aziDOVGZVyFcy5Uh12h/0vJbTfWOrMsL3ZsdjtUXt35xCNea5JKB3GfiEIJ/TYmzZSf
YhROpA017CshizAMNEKtAAI2+Bdu4b05NUYWg5EZoidU6EFZI1vv0oyOpXOxIT0pBHUzvyulksAO
ZaSzeUf3mWFqf9TJa8XqK1AQviKigrxNoBNL50AmFyMCXQs55HQNzg0gHiNL0kNLc96Pu7FMRLfX
Euh495nnO6qNGFBXcjGk4LLu746R79UcrLtKp/PWf0PdcxBp1TX5q1D7oQVbZjY1O1ldzHyOAQJl
V+ycMqWZqO2YGZrTPZhvF1PqjD9NM3L0zv6RqAqHPjjR3Do0Jcro3k4nmt+D1zfCoCC8Bgnycjtz
8wdsX3ZyKtVEp+n4BOq6jY7p8Tcty8DxVJ5CaJb5C6wcvTbZgCse8uGBY1i6eZXnMdFAcHC532sI
/m4J2d93AsHnU3EA6cFclBowecgoj7gfUmOFbemgdEebyMwusnGEAROlPMEk572gDhL5cWADraGJ
SCfBNwS54VPePxVpNz8OHx+n/P84rt5bbW/TP8S/XbtthJaXutRKAhAgBWFsbshpawF9OqghiI0U
V2AGCUp42ij4femMOgCWETi3jy7ceQKzfcHjF8hbmILIieN7QvCHaUowOr6ML4RxMKhfdiF2gsfH
Np5nyis4407X1+6T9MeklxEk8d5vBxYwxVUdnG7uhkDUDkfwqGUYrwmaBGdNg28XMFSSa1j62Zzk
2SgWfseE/7M4YjNtccG5YffbQuvYtL5BQfN6UWgi+84sV+7pL6X6DASdVvD8ZMxIdtoYDLf0M+vG
KWbECjv/f4v1gcn8uhkMduUdB5J5f4/pYGvaV5JdaYXnxb7zF1zf0Ge10tPM9lGSTugTVNH8EXoQ
zIkx9LOnaVHGqCCp0SOxx7pt5gvycB4njcjnDcNE1/XEhEyQa2lIn0JO2MX3A2SbdeWrjvNo5Z6M
eaEG73FMDp0zW6PEGSk4lM8px+RiM2P68+wehBncDG9kgBMMIrTaY7pMO4NTAckOxljoUfT0kdii
4vNpzn2wfcsn6m+Ag+6H6NKBiXQ05Vs2Uzbhd2RmEmP4RKP6AuFfLPvLJLtNIANwQmm/bIQXMuCs
26VLbzduq4hetiRyyzv1T+3jJ1dNsAk5lJWIBWwW3qBe6wqedP1pzU2vafGBgnGxboAmqv5YViER
hlJG5RX5I2mInoY8CtK7ENpqFp3ai0VL3+vPbVRn8v9LSOzPTGti4CUyXqxbCIXYsbn0TqWKqwWa
nEqIy0RDDZlGPzQytLSmRnEGymPUj5C2TkjTOkXR6O3YJAM61E4ZniZRS32YC1xhARZAdmEVgc3e
AU3//IiToayJTKhwYWf6ETSVQHYHu3HRNlsA6kT3lUDHeeL5eB6AIWfTD3n7XES0Q2a9slvS7gdQ
QYMcE+q/rY6q/yPdLnvXiKyd4c09AAbGsaH2t8c140xriGEvcUjTe08BoxKU930OFkduwtkys41l
Jonssg+o0+tQ7agnErD07x9GTbGWGCy93ISXjambAOChmf+x5izB+kGUJllu2iwF6YmwfNWo2vY1
rHA8nlv5X5chh+HgANvT/DyTIFtysW+P3lV2c5aAIS6SE+iqV7JUDG8rnJDlbx2DMW3Z9K+DVn2f
NJYEpXaHMDjP9CiADi2+V+lJho5QeVdyVY1dc+jvhD0Upz70MIti2uyUPjMZZFEYRXioU+w7UHBv
ou94C2Aw7/B0qpRKlNxWW5JPkUi0LjMtxr6e7tQrmSdGhrTDBXc8LaVHZwp/dn3yPp/3OL4T4FLB
8U4JB1VlGY9bdM7G3rnrMKdpVTt/poVj34PJIO75TqMUvct14uwKx2jOhAd239MegkFzt//qlHpq
qakshQGELggfCixGZ42lSii0S8thzQTwDOOUlXkWS4JPaxt2bUJWC6ssikMczV2geqwnUI3u3ron
yx4SvUBtlvoJ2o/lpPqCcaeDH1KgsiOdxgj6x97tl9tgxyWpg5z7eW3zoVZ8BAviTXFBrrc6m2iV
QLETYhcdEWJI4rqVLQDFBwawkIgCaS5rC6rfGGysnnlp7pasDJyg3zi5ZGf7N6XpLNQkSNw6Xcc6
oxPEEzC/FHHBEfQKfTECUzQgGvkSx8Kx0sdh7m2S6GvqSNKGzex3nuqiB1NvDL8c/iPbE5E96adK
cgcacoY6NXGA7aTIIEIkcl4nPVBq/aL3SV5A5tk+ZepZ4P9lWNTIcPLP4NVAH2FtdvwSnfu04kEZ
JVUagMHb9js6awK8x4MX8Jql8uFfHNgNjw3Ub9Btk1t4oEe3caEsUxLcjpaOC4eJlAPBDyaPc85a
OczBRBbzDAYu8Xsu9Mry3jVtbM/zDwslwd7wrlmUmsya0WM1FiaabdjxlBNNR2S29Wg3vAMF6BlC
SzeNGDUTOSSGwX8d0UIY+rs5MPaZ6iO68XSbgw6gUbGEOkPafzKMzvW85aGjNimq5hvrFCpAoSQ+
B61L5jQ8n11qTZD7sgC3oJ/l05MK18shWBn8TDZ7ijfVfzSfyWlwfWem/lL+Lijm3l2pTvHqM+d3
UszEjcKQPzx5gQTOp/L0b+isnXRUN5DsoqRDyIuDjPISHObILKf/+UvUGhAkF7nvpy2B9qE1xsZM
PQqJW/8iiVGrjrZ5Zm+N/RusSl9WlIUA9ijCGoXauopSddYwdLFCh8n65/ph1Gj5331+e0a7j+mL
66MRkCo3I2OFOcTOXlmVtvjVOdB+Ljh/WJFwlVRdKLhPvJ962C3wzAmZ6i/R9YzidOFw+BBHecKc
fb7ZfVeMYf0t99aVRICkTyZ5z7td0gEYHIyo3GQsJK3JirWwtyCBFEiz7wpRd7dMj0GflqgMXjnH
cs2bX3BDb/o7NvHQmh7B7uK7hOt8+vIU3kObT3FzlFikU/ofBWHhltFe8HRdeXn5/FiQFlSX2TYi
yOpiJ/yQnbh4qNwxC6X2FjdGx4smg1s39rFPgg0XuoeG6sMC620cOEO+309HiMQlapjqhsf8Q2zP
GhNnbSmn+TQCmLZSX06gD7dl15oSXJ43dHpqRlbHLynUzjP7BqZl6PePUIQ9nIQDsK3znzXe4rxc
lNvSeAhXFI9uCZZtcim/sW8B+R3VOW2PX2rRpVXyM5ZUac3RA8I4Jet0uLf04lyV+ff6Vbe0vuea
8/lzfimsfu56rtRc0s0ceGc59LipydnHw7PCOlgerkX6dB4bvAH1IGvrDVM1LV5IkDoxjszYQgsJ
3Zgx6APQh1Q80jB7HqSXbdmcrSLqe26clykfGJLyMgQhOOcdqsHBemkUHyVt37YTIofPk6wWrYpp
YNnTqRKbkLDUsfeyhVivW5yn2pU1vn0NNZTxWF17nB6DmEmY9LrCRbDu/fI7FRCmKVpTh5m97hyP
WAjy5ztpzcIaTv/VpbefajwH5vxEUPsRA4lpm2gLX/nltZCPfnYG+vQuflQoo4PM+rmXNKwe2/S/
svW5tLykaiwaukuW72x+KCGQqWnK3EH9ZgvMbdJsULjDviFKJwFRwrp/RcD/AeBXXKSpawHTD5mR
L4h3hds05efJXUni9r7QqEodjSQNlTQ2+pHc0tPDPEyU3MWXCapuQdZVqiBl6UR4JIC+6eGIkFI2
f8zAZfYKJwi/2WV6QkV7CP3qN2yBVB47s1gTt9LZFJfpZyYydQZhg30jqFfRHylnf/jKbLbxxMIk
mxAq8ItAteJPL9/rKP8u+B9UqvEC0WaKph7u8qMkujrlcmGP+mOmaD63coEDhjygX9wFBZK+NrW6
Qws9vgkAE2fEVW2QfcuQlRbH5T4Rn8Lxv5gP0jGkekock2Zj9EDHr6RYZ46eXdgkg6IEvVnn1cNF
VHcXa7670Jy5OcLoyqHERpMSYZulHH5kzBiVRXUoLuuG4/qsmfSsYglOuqO34fDNBqPmGjF5Txv4
5b3eAEHvNitGIY4LYDc6Qllz9nCUtEFzJeOmxS+8NTwq7VrIbEuSPdqGN9Uc0noGu7xJ2s1t9Nyo
S1Itk0AThcNH4MW5NKLfaE/ms+HzZwWMlwQZn4xzNIR+XNWfnKKXrRnyUSR4235vl5hihkfuvM5l
uGe218spLUQ3/+SHqPCemWh99fIkzISdC5UQYrdw7XR+kx5PEsRpK8/eKaEiQraa0kCzfZk3afjD
q1KX5Zgdopqm3v0pwOTy+2mQ7aPhRmkXzo6rE65P34+4+i8HauLU3QIViqY2nMnlFPe8WzJEqkdT
oycj6SenXUXoTXdsjqHgIJBR3QSg1AMgqI5LY7qL3S9KkYK/dbzpt64xplu4mWf9iaGCPDjyhhh8
IRIDRKZVYshIGPI1Fkc8hjQ0do3++2g+7Gpt8MQvpewSLSVuZapA2MoWwkDNcYs4ssIWOfUIqukB
igUmuSxL9ioqONHWcQJAkN8DifwR9rCXz6fOmrOQR/DijFPA+QWQaxn8rS9wzupOCfKoFSJpjvfB
K81dps0Yj75cLpLQXHQYST42yhyLuVAhIrwZ7ki2+kcBUnOsI/RDy79PzLHNAEvQBb84ByweGZ3+
if0wZAPRjCaE7HZlojevY3ppV4qm+RACLRV4zWSFwn8pAKKa4T9g1DiXjonpSpg7zl5+WgwnCLua
ThIf1ya+7Queye3ITjooBQ7ZnEdeSRqwtE3lUsIH2i0kJTs+jFdf6jAjAX8B1QZbNgRKoMSUTXea
HpIAM6V5SN6w0Zm6ABnXnBeyCjxYERq/LDuLCVELRv2CX6NFDS+q8Q6gyQtiYVqFnYCwEXuYfHXT
hZR6dmDHnwSADoRmbD/K2GJ1p53WaqZ6kicLwOJ1TsTXDj87Ol9Crh6u9tmN1mRM+e6ZngLu/1bY
drO4f0uvCdAAqWLq2x9lnisIkjFYzMNWj5/ThofAw0tMZmSofKf3ZPxZINlJ0jGpqjuo/fMOXVHl
03KGYWLIkTAi7cX1fmPiqb60U7fArQR1aKpPbWl/DhcoG3cMJcqcuZb9Zohf5FF8IZUSpkLvKUfM
fwmWkLH74Xe8NUcjBz3aehQ3bJ7/U2Ywq2PUOgnDdwtlYzJoB/puSMoHFARgGq3+1dRo/t1pUisZ
isLyvKJxcL5eWEp0e+khihTQ399G6R/NTebx1eCHLAqoNPItJnUA8vaI4GbdCVITAYeSTwGUsjmg
qh9ZAlmYg+vQuUF0zEhY5JjkyvdsCo1cOHQ1yMS0Kh3Iu3LQKsB4fIwyLZCaFRNoy2dbuOD4c+L4
HpqLYbYbklTyGtT8d1hW+Kown0Yco6zebbm/fXw0jNV5w+500PpiVQsKy7RFn/g37p+xY0lErYo2
z39jbqax8yf4tEy8i+795QjaP36+/eTnDqs/GjeXYTMsacnei3qQM4oioRejY8TxiNqMqHvjCzFL
0AllfVmPtZ2dlWwU384QtCwu0NebE2d6vDODD01yGRWDFswnod2ur2Wna2a1KOUjM0/jm5aCR51G
9fnfMdtYR8wnw/BV9vwinRK8+iufD576nxytqcUQWWHWy9JOFRoaBGmF0S0kuEy/0XUujSmyk2Cl
gQgc3IV5eUpv4IE9OrJXZV0rk1/EAUngjYRCcD5O1uPyvXngmeJfuKfS8zzm+PGKc32NhZhv1AiA
Qz17Cf2//qAGQ77r95uxdleucyihQSL0hVXZcVTY2K0Pe4BXx9pLH08kGfqkGg8pU3ti/u5Px7aF
QP7fvuCoPti6dd5hRoW/mH+c0uXXM8GY3bKF9oXoC/gLzLXwVSuUE3YG8Ef7KlCQfituYRxN5Ey/
ggYUoqmukTbTmwl/DL0IAQ5CVtGDc4DshWuCUBrk/gQimEekQ4OTzPYTSNyGK+EH40bg5j5gJjP5
Yaa9Ql2aTSHRDr6gbyES3i9d22/sOZsvscgbWGE6LkfcxdYpxbt0WQP88wLMeyNLVub++b16Pr08
qJtdrkKvcX67dp1GEiKcP/tB0KKG9lVw1xuVcLZPWq3lv8Z14XGs9uwLvvO+SvKmpDbXQJJ7xZJ1
QRoBvLfW+dmf5PDg+SoWPrh9a56MHx+0eRjTrpIs9dd5KHww67Vg0BKR6U9cWDadZd5uDm6YWnk1
nwBGZZ1n58JvgJX4rYIC/SnWpRDxjYYiwY+ZGzrVeQUIf8ps3WP4kMTRCWcgEp1hz7HvcZXBk5gt
fFVDtY0ltkUDQ7SC+hXcXlQMFJr7/rgMSee3oMtfHUhDAZ/8jzxmJds3HyGjb90cHFifjq0q70HP
HwGmyR1+faQ6ML8ww6BW8aIDApQmI6R+osf8oxdqWBRHATkcV7GEOb2B7OSsK7Rs7TWbH2fntdIy
DKEZpVHM2IXcvae11aGRxT86aRXua9J+czMlxzK5GfqsIbH4qQvbjAfFSJnPxvfqiMD3s7bMA2he
H+VbOKDt2h1wXJctdkgg+As6YdHhoxO/363kjO5CpfwixaaalO9sT0Szb5EhDfSdSDgtrGy/LIc=
`pragma protect end_protected
