`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Jo0GTP48lurGV9QI1c62RTUP1YVEamMz1VZFzIOsgfj+B/Me/Uz/+TNhvOgX00Boh3rVDWY3miWC
6dvD9WUK3Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LQaetkHlTEQ/O2QuW4ImDf/K0WBzrX60Y2eOh0Fzlit7V6+gYpu/pdjpcV2iUJ0OSkPSJI+Mhtnw
My00nmvcw7hr27JQMftgpSq2KJTPiuvMTKQgaTjH7G11dDQzZg5OIfVuhiEdrvLjBL6ODFpLjnot
+wtza061w0h0SULGF8g=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e7yz9u7SkKHpUf45ToebPKpSB+7SYjKyIPDWMVo4RpE1fApRY5i+m6AdkyczFN3egPL9yuxMUBQi
B3fcWe1KL481lABpqgSqODHUHO2V3VOpcYtVbs+ITdbbKzYLqgggxX2OFaFxfaKpm8KQDKkYwb5s
hDH0bmxkegiSbK8/6cCO7THsM2QEi5MCtiINLnSFKZxzW2n5D4XuM/reG5kcwrmcvNmgwL09iDms
zsLNFk+KlTwGLQ+sjNp4XMp3wRVy8au+yG/ZaAjv1SaonTr0s0Ktoq7kpKzzK8Vdx3gxl98oC7lG
qI6lKENHTJsj2Et1sJqARwUVTfXhIwUnx7z+eQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YUgiCLqe/j/NhPlORdPixdVwbLBtEL3BY6gCgf7tGi15P5FTCSoEIKV1fMOt5n55kUiULz6ixyOx
w6KSNkCTxNK1tRyjWlYPNwh+30X1DX2lqxQedujI8dEfW4TThaFzjbr5VzZ5Xx3QklpDtemVWlfc
v+85sRR7dpK2+yz7JHTpwsBUmUIz/yQuKTPH3TXkcTEtK3SDtuMd9W57I7EJRQs/QWb0HRC1gqri
b73Bznz/ITOHvk6hyVhz2IcLVxpPIWw2SPni76CtRBGxpvEkYBsB4Tb29iojsozDmdeCBCdMwy/R
z6g42MtTw4HdwvXecIHU1Ps+g//YLogOmAG9jA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
m7rYtXUavsevrUPbAA9ErlXCOGGk4fAoeRrucNOvvuTkTuigciZtMDGFuNCCP84AUenq7yf+knfr
YxGJdpaWbSksXpHqc2OaU9JxiGbOYXsVLB6aaIcsBViJ1Iu9Y3dsxqVRuEf/+KOaUoj9MgYpzlBd
dGJCSN02BKWDuiELCvkTzxH0HkaQw6L4Fs4eaqtvZO6JC37ps+GYsLvCsUVOUrxP3ZXffR/5rO+/
r+Y7T74S//4yP9CGXNTnVBNea7FKmyEzggzbDLVXfwg7DC9jqBdVLhJdArtJhH0AWfbyCLDAfF69
TIFn/nOkcwqHGmFmfhdLuMOHq1GabkUC03gqCw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WkzTVLle3kbJDg7jpvQ16rMwFjgKsN6s5VraGMgY5PuWLmuM4CseW8hGJcsf4WjZloefR1XKRkv+
EV0MnXlsj7dM99Z1mYpSYEt+FSSlVw8ZrTFDfAXM2tVaQ6tHWq2thbcjDszMiCZNwxeaVwffojNF
dPRWtPW7gJ6hRMZJ1oE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nB0LvvHetoBgxBsMSEPN44HAKokSVtsq+whVeE4wsASFbqJ8K82xM3hbmxu6ZDYkwRj1/AOA3HVk
G4ilfKGLy/G7TDbQDfRO+5Y01cbhrcP/GMxbBzv8olyMaD/JTd0uTncjO8AIV8tUE18Kj9ZhfRCb
zatytXSeRs9JZ1gbnMMyuS9DWHly6IquSzk4ICOoWWjyjXwHRFPGPkYHKeAKIXuBgNn5YIUb73Bg
ZfSxBEDnDG4lR9r5BsXVWXPmkRPzzmalgCEOM4dNamRFXJG6Z063apEzsaFADjlPswBxcO39daPt
PO0nWMUFnDtLtq5NhL5JcY8vaGgEnfVUj0929g==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kx2/4FUG+WgpOeMb3Rbb/cih1lc163wBQ4vKkckklmR615Brrk0uvh47GWx5YPIQIJ1dUYGfGof0
suWssmlsLprBF4iyZ0oJN+doxvhmSoNuyqNtF4sOBh2mA2fEVAiuuRzdRQMw/lsxuNxU5tTeu4Hq
m6fseqlUS4i/DqAjB6NT+vlMZPYsrIaV5xH4A+ZthsSp/Yv1VhT2z1Yf0I1zXIDSJLePBat4WiXu
ztJa66W8SRYkuIFjEUecZElA0JE2MfS3tIGvepvw+Jw2NqcpRNOyHazWtDF1qGPoplQ2+iAwhvFE
swC4IvCafgzOO12FbZwI5Wi1IC0+7hrnR+7e/A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135968)
`pragma protect data_block
8GvLC41uBcFwr5Ki5OvQAwh2MwnGKfuE0FkJhaohC6KDT4SH9pKcwnvFqbHTm7H+kxpfjlg3NYlo
R8dPW4XArskiR6Di2uUoB/KHQZgA9Q0cwOvSEJCPXUoGkiXhdEHBdZvay46oLEJfDZyIiG3DmZ7j
QdPLJCS+XMM61IeiXEl/KfRAoZPcBaiT0WAOfjgCAlQMalNjg2+HkNE4qdrQ5iqZR9xgV0C13qvm
4XNo9wimNjkc6iVn8etC7CbC7MWQ8oupMWQcQfHfK0x5Y13QuMd50gURQS+t6B/q5MJ1P4JlC30X
z90SN6VpYl+JjRGApMdhLG2XqG2OQqiExOLELqqXZX3/XI7gdW9RmCNsVhZI1ervByMpWiQPqcu5
dcMdsX3Rwfhr42f/Up4DHKbIhNhmS640lE6Av/wC1p0PDlYR/DcEgwsVvG792/L/kjWARfhTLFNW
a+6B/F9fbZ8gmm6lHquYy4/QoErvdDezkTtX7DV1u+aJy8CR/dNR/cnV9atKRihc8FwU2UK2CMUu
hSBBW8dqXSMYoBweRdQ1d4EjSOijAX0hzrhrax5VivNSIBlMaLAyskYX2Hw/7mH8S+thkCKPD1Wx
QSOHO65bUF5W5Gj9jSnPaXTWgoqCCRNrnO8tRk2M0JFvZFb1JpEVrGWUhuTlnh2qKIEfUAHYEqjQ
WCNH9tgSVSh9p2I8gq/FtbPkS5bCEby2vSVYkS46BGo4XvCrev5c0HTYD4hAB8y8Dc+nDMoibtUu
/1cVksL+t7vOCVbtQVXLasULSIU5GGOfqHM2C5tcMtNwrOaXjhXs8uGOu30gpf/HQ+FGn0ee3DuW
8O8pAMKpUFrwE5lcgo5JAXquJWHRQPGmvZxndIib/h/gD1RJk8lFZJNe2figE5CkTc3b4gitsjpC
qhFWBE60g4lRbGISC+cYTh2ZUdzk2qceT6w2EauxWNovCUM4NnhrHLb98Wly7bngvYsJfK+xeq8J
qd6olEt+T4CAHYJECBRUbU6FBnL47mwTv2vaAOsPs121TWNT2ZlDSE7t2WGgORH/HlibFgcm/YeO
ddBvMNowlV/v8QrzbrMaJDjIW5Z2wdJzUJH5nbKF+hPGoAOFmMywGk3OFk2lYQ6NWUPoBVbdeZhS
sq1ogeiiLcU16NBofhCMrZNqnV/YfLAPOWQZUUrmovHgTv/cW2W6+a132IIeIRCWOdvGUkZynDya
57PtShvHmZZvY2zTi6c6OG6YjV6OVbwbUPvAY3gl+gsRuQyKY3RuLO1Cqe9bEhQR5sRziEuFLe3f
F8mVDKsnbFP+MPptqe8AlZZF2m0fkYj9/pkc8DNpT+WViBlvEaVGXkSXyMFA0Fuk9SW3ata4eEZy
awxCaHa+uPkxJFlD3HD0LLsJSQ1WwLh1DX6PtmURDHeQYooYnNBQL2AaT7N/7xEdayV1j7FboR04
/KStsSkj9nQc2dmJeXM7UyAkm4p2ad0XAyFxzeUv1ITQUwZSiDaRg+Pc9/sAvMpzyZD3jP89yeoE
9N2/dE2daaZfEhCGtzsmOcZolrIZCsAMz94h4CdSsxO/qfzWqlNgVAtmm9/Fuo9MpsYCVWa3HzGV
ZMyp/Xe+q1Vpqon1/likjn7gJN+v7rEcXjqSr880l4JeFfj7WSLPq7Q239pFk42PZxAQwzWmtFGG
Ky1PxsjJiVwwpAuSvh9CYD+LB6zi2rMIOUyAJfdEnl0STn/CGOPR0ckyHVKjBN7ieT5+z0hBMr/N
MPuEyHAHSfsbjkU8Dn/Ypk3IvEPDTOHMYXuq1k+vcQrXFQrJU7X4M3L0WQRpT8c5dexIunBTfk0d
nWyPkUaPGjJmaJhJYQ13JrKKqsyPxEOCjK7xdnzf+ukNDsf4m65Z1ATXa9pIgfjNZdRp2neKkfr5
XPeXUmVrGGozHu3S1iIvAssyzpiJtc25+uEdB9D/IlYmuAt1YTkXrNprKy/DJ4bb643s6RXizLg5
Ws2lVAgLipT3n5sbEd9ZUdaPF0mn0sD8DIath8vTfm4qqrl0Bk9Cei9BMms6iXLHv8MFIgnpZ1Fa
ZquFyceIp8Bba5Agz6t+vUYJwnfRbqNFhwl450MxxCb7Q60MhwXOzAp6gaGHpyK36Wxu50C1pSaE
d1fAQj7C80OCqbrRKJ15dtp284PlmBECwKTKxLC1UFD+49ltBxOPWwwjik8Br7W5Y/ZvcaAqPNHM
ysmPkzN+KU9zWLWz8uwOrdTOTzJBrm2FC6eFRl6MqRXYx2vNw8FHBF01RMB9O6UOM65CRRFnmDoq
2YwrCirqTcWlGHBDIk2pNzCQ2rsmJ+EdTNCjkK6G9wm9pS8fFWwtugBQUK31dANI6ock2i38+aoe
3smZRdUJa/dTX4xpGQ04vfl1EXnuxK7XaRvrf7RDiqRxaRJwVhG1/o3daDA3TONZhnRFbEsQ7RDF
xCJryhDwQjCWHmuFfz/HcUVhGEhFiCjZ1K/H2JbxrRreXBu9RtJ5jj9tmjaak8W6Si5l4WwWzhJ+
DHOxVaAvAq5qvxKgWP4YasDJgI9JsZagk8RKkDnVVM2xzewfFvnEqN5tpxCzXCBfGxE2AdBiioUP
dS+c3tASkDUpZfmBPA1LQLeTlU/1Z7LaX6uzERoiAzMZQ1x0u5xw+xxPW2m6kg89Om496VdEuzg9
FCTXva4D5IeXfH6c3N+KJIlDxII4VQtfm8gfeWAdRhv6h1qoArVRxsQQpKG2cjWnZJopBgW2wS87
dyC0KF1/dttEZi/0h6X2tDJHDJd+j5B4ss2M/fLqQoh/wc+RxmmrGqwXXCxrxSmsHkxoxRHn2hvx
yC0rTNMyvwfLDfyqFMKBxPLs4lDaJA7D37JpjmsudRTbhChLJtfGi6OziPDDlTH1AItoakvxmhAP
swboaNpbPW+rD9e8/2r4G9mUWyb8mTJEw+puV1ZS3fVz/ZJ51GA8DAJLY9ubfNWj99ih8xZfMcfQ
NvMKiNw+Tf3Z6rZtFy8OB0CN3oMgobQVuxib5B4RBXzJAWfmWM0aUHSTa557UdzGl79sR/9PR7XH
4k3bVAYJ+GWMyKkZfNgPYA/tepEzFpHqtLPCSMrvw0/rjMjOGLRFPzztmP1Zs9AFvLPct5tsaU2h
KNaJghxHoLFPd6gyP3O18/GJeCuWw0h8RmgTbJgcglc0gVnJme3xhqI65o9TWw2RZCOEUZ729PV7
1H3ffoI6aQB4TTKGv9mVuoIjxtlLphlw8smvLs1QK2GzCuzh2vrHUwvkR9do8QWmjX/0j/Mh++Hf
4li0JMAwdkRCakCMsLp/UDDRPbfTeeZ5JcBkNO4ZIoezwCMSztanhnoY08uVeRzGblRP9N89YIqB
oAOhwOqDOHKbS8bDvSgdMBFgmEhPlqWyDRcWJRxaQJ669zJcDMIjZQB1FiN1ZBWm0NPjheGEV850
fjfA6L0y1lHWeK1b4CD009novv7oVGFmrVqZCWYxd/KvMPMZLJxNmBB57eju2h4JxCZqNxa5e/uZ
vQ40GsvqOgWaMQCM6H6pVL7fRmXN4PprGINMI9fQAJbS6WuXTXXxJTGYdZCjJu+b1IZwr2QzHBSL
Cxy87Yi7DNrtewt4AIpjhXiL9U7ldVBDkf1Cf56kVih6ApRncYsDD6BrpqsjU+diYGekdSXc/+JH
IAfaQX0E7d+dGELuJ5K7Y4mf2GLmtt8XloP7GC+cn3WfWzNIK1TotXfVU+KDg55Fc96xnOuS0CNW
stxsjRJuHKyfzpM/GVWDxeqp0MCdRWEPadDlR6FlNX7plgof4A4+w+X1CNfwJZuv+c0DjWPUt4ad
XKn0vZ0C92BO4cK9tqk6HxbOlHNipjgeGyv29S7lhiyhmqRqd8VmK06pr6GP/Ey2rluIisSBoZGX
7OcP5qERSVnSHZg9kHiFB3+cgw7dCCQLE0eGA2ilJCelfu5ikF8ctWV3mTPCIUWapVTLyS1tlohD
pN3LESdL3U87I532VQNJwPuAm6WNnjLyn24AxqtDFW7HBLtrKA41lzmrPz2jl/I5wffSOrUmEjMv
uz5m22gRPoQQ5noVO+/Roz12f2xwyNVq/bJ/WmzA8WZuCpWXDVfmm39uemDUPDlIA7rXD9AIS/L8
O/A1xPqBM67jr3ARuLIswO7wBrv8nGQWVTh9Q6go6lHl1uKXmzJWHcG0eKnkfGpszdiQrwuGjq/0
TL8IpH83H/3c1VOAT/4AQ9FbFEEPUblPu1hAvP2U/mzO3B53mpEae0y+NlLrBwD9WwDrkFtfDUN0
2a8Has7fENfgBh0mK5+7BMt0Edr8CQ102OKJ/53VI6nIuEgyKX32J69KnFXdaUbRB8w15oznZrtZ
R+ByKT8R0jHOFIajasOImiuyZpYE+pobgzTo7KQOWLRZ9PhmsvDWN9yyIESGZDFhRwQShw+WBrEM
RSp8NrmRhHBp+lWfGU1J/4J7hHJz7nMBxaYy3n3XD4K9bF4Ymar804QsIJFhPYUD+sYrxfvh+jqF
6tpOoYhPvQrnBnrTU40yhd0dYGVqVExRDEjvnyIV6ta7+6xVGOiuo3g202HueZ9iy360ED7tgDDT
mPM8g7GaxOkSUVoP3dGIUeOXdGUPZCdsAu++kg+wfe7cGTqBGqXbl+oZJsyfwF47kKQGctRcrERP
gE6rIA7sb9R5j30UGS184yqkPayMXza6RIzaGYdCyZMOZ8hkxnMHms2z91HVXhqwxXN+eBgKan+s
d6BJXxWKkBjvT3EX+7XeRH2Fp3mXB7f3TqalccHUQfWUPOxFfauFOsFTiPQt3cwR0UbPdXf9Wo1f
wbnBvIHER0Fd7I33vfU864Ao08e5JbajjY84Syhp4j/IS+0/Piz+4x699m3DO3aci/f7hLXgcqJx
BUaDNyspe20wQmErfNuWONr3twRgV8PiRwNxX0TQIMHFypYn0MwC4IFX9QwwTtSQ0uUuYwmPnPib
4oBFvQFLxwdnu6yI/3j8gjH3rGAdIsSZ/sFQm4EJurf/hGAz8CuwdzhJWFwtf0R7SQqjxSSKbj5o
Q+HJ+LmjPAgjtDqQ1HmCFdTZbQ8yLKilqOEPfxfoF5YDIW3A/iVRdWoH/AjUrcL7kWqtAe0wKHwX
YdrMgWeO1Kxna+2JMXfMmeze7WzBAgSmC/kQ0ZHZwmS9421YlUWeVR7M9vKTPAcTMLMjUV+dBIh+
S1u+4eF4Yb9e5virqatBsp1JpMAnwXZTvcupN5Uz23IZanzcyO4t8oQHYVmZk8kF8ZdDJk5F/PXH
Xq+D0sGFTiGu8z49pY5S/dUGedSjcH00W0PQVzUwyXVBXB7jWmbClg5bpdu6N0tF3bbiRiCLa2yY
qVmwhwG/+BUGyHHgAKnwrwPWSTUXRKsTSkeaIq25DB8B6JypFtwhbUFuEog56+eyNZ9BAeZN1y/p
SH2BGOQ+hC8pZArN+Xn2Yt5iuHKeNoftIFhHCwI6WIHkzC3HLhnGLib9/ghoF5S1M6+gXoLdlV0I
z50TvFbWWQ161E7zbE5HK73eWbRtp3Ok4Q9dHgML1M5HPN7fVnqokG3HkBLzoTUOJvFSOeng52My
Js/CgfskSsVu0tbvEicXxlRw/OFInJ5qqD+8/cVICuAZe0y0of5pxHGoGAW/aJFXwwWjaMzCWxzk
Dgl4PtJGDSMQTquEd23YbE746HVdDE2dqI2n8oR9OuF4vs4HjNdLTBN/rnUfu+QJjGpqcKE6AhHb
rqltxyYScS+3k3vzkudci/twcuiJCtAT8/isuxpuS+rCfWIMJjQhv3aMHZt4JC10Zsq9/O/ksfbB
vljjVoyeTA3CJoxkjhx4F/vf8+DZaYhWz1uR5UX25mPJLxZ+vAUv8B642WRnKqpWQBIsei4PbQM9
lioPnDBBYhSJrMEJj5jI0A/n6vdJnMNEmA/DM57K4oe92awRp8HDdA0OauZrHSKCeMfNS8jG3Y13
1QXIfR46rQlZQng8N2hNHIhUODvTQ/d3Pye03FBvjGuM+uYHgAzLh3PIUOLK6G7dTSaPWBTU3aPU
szo9VqJTvITEHbGvLu7NVJKoP+GxaFmsSKCy9DVVbYRaMVwRATt2K5CSzGgpmTdhiGrGxVQ8ZQgU
7u70Ly5KEW5dgnmmswV77Qde5py2vE0gaAjdD7m9QGMfAOvq0E5glSmH9ASb+jRtEBSVX2kp05vl
+8+N3ke+9SGnGHu8ZaeSs1Ow5npRF/f9ND8Jnwlic0ZK328LVIHSGFqQJ8u8nDkE4M1CKN5VE+Ty
n0xEI8Zk9tBcIPK4sf8fD5g4NfhHT8B+fzI74MWRP0fJ30io1bzbGT8k9/8uoJ67IJCCOfpOkAqQ
vMY7l7wB9RnBGx4POUz1L819tuek0y81IPNWEYulq+bURb/z3YTzZ69GZYTHGf6VuyPVZP5AhJKK
qvXNHzrWm3yRYE1F+Qju9HN3is789fbD+MvuFoWfpta6Zu38C4UW9yPXXz1V91wvEYZ5nC3QWy7K
ZPHRaqkwFY+kNAQLNR/m1/TcA57b/G0bZrka+pL2fX9jlcSf3nbCaa0TiUR2gMGHemN7f9AaB5sc
8mQpL1afysYGzeB7hGDuwH6tTh0Le7virlT9UhATewVsxQGN2Phm9YXFJAzMbH2IPuir8PvAQlxa
0x+wkQ+VGxws6TR4W6n5degEa5ZwCCKCMlxF98bd3REM2pxRtDdesRO9x7Z4sigkmdG/esTSXdLx
J+ILJ0oDQxIiOTUGt4TF+pnxeabszw1npXfkpho909lN4+JUUaYYDc+mUHgmEcUeqQkE/kFfI6RF
Of035I6DeH0HI78GhvvZO1hSDCRfHVzfksoPDjuaqrIM7N1Wlv8VKybzN8PTUGGli7WP5NTjrVL4
3wAFCDrTLoNE+iybUx7DsZ6/IKjAC0bQu0aWqu8ZZaZlfiTcbW8SpRvIoIflIFlBmnf8OVFOD0Hn
CXHzbuwxRprFlQIp85J4OUDmfkLtHRp3eYsBgjVM1NytXiEsauqfWucpYRdNxSFYWxFedIl8F1ob
v/pWIMAshNZmFhg82Tz41VoGDq3JIkvG2Rf05AaY2+jSeNMKJa1KbBE69Q0R+/At7wylHSqemuG4
lFZC+kEmG3qqnt0HHWOoFB/Df77NvFi7rXmY3Rq/xkFd0To2iu5O7ZfFdkbkzUatAeRrVBqaDdfR
hPrizQYG+VzJ9I6kVXWAQdMPhzAmU3AL9ek42IYmt02Ho0JdmHa/CFLLAyO9NydwAGiTlrI25gtf
+XnrJPgHf1fpBo2XKjFhtgR/XYUKfopVWvxLrLAiTAxl1QuARsYx8dst6FxMRIHJ4eBorjfGbypj
rDr3elYYm5sPXAiZ7XbkcpKFLeCBCEqUwZkMeB1RHmeOm/q6z7Eg8+E8TXgQ04zw089s2IsoBONc
L1sgbiV3bNXeuUYQhKt1aDFcZYLVaQN83wB9Rav0iNJrfa9A+h9XN4C/Xp5ABZcHesMkJ2BUQ/N8
LrmyeJGJtNncVeoKv5ZTzsknfdnJGGzmkFdHVha2OLxDmgUOXVEb9NrZq/yAxQMYLEbaqTDtVS7N
muTK0wCs0sbQ0nQgwfzadsxKo8PI8QGCfl+L32cp//HMYUBycmZwQONjSLTzY7weOjhbf9QtbdhB
24hmrUEHnExRKrMGJ8Oi8fT5k/c//cYw/h78y955TGWyfO5FYpmOLfs1rzIceYQEmrsHAjgLmqb7
QfNVDpjVQswPpgm+dc4Ckr3LglPEr+D0u+z22ToM3/PcM3cLgFpCYQNN4zE9q8/jH3cFszoNyOUZ
cQ3479jOpUUrQ2Ejvi0KjP9yQjhwGBmjJ4QVq0DjNmTiWYGKwVg3UFoUVnIiPkcArYgDdpQhaUFR
ESS/hqbY+unbuqNuJyI74858YFfFrNLKoyNCW61i4Yy4fgFvKcjUX0brx28TkdZYeOphGvJ65SjL
mwNKRWCmGGDHv9KZPxpEoWs4fhWK1vmzs89HdYcl9uXm/bG5XP4OgC3PldYOgZHPLiXL16G+OU9n
LiB5BkDsmiDUIByKgi8aYGKflrj/gnM2UtRmxABVyadx88bpl9HD2X8CDDXL/3C1W02jTnMNtyuy
y2vApoKE6QjVkW8OrxJse+xQtCpjsgRbmR3zdsxdqdsEUFtW69IpjGls3W7glbm8j9SnPsHWwKHk
Ees+qad6kDm7yH8k0XenrRwLI4ktdjwiJh5z81vus5Zw1Xrzed1H4UZL3QBy7/Nq9xMa46TrQjXa
cpDg8+LyspCPHtDcL+w2fW+t9qtYwxxj61wVY3EsQo5o/yWJc44Mbx/BJsJ0rFA/eJfB25xEzQey
oMLjnu/+pboTWVkk9WxdAQ8cEHAM0cRkWlFJ6KFDrVfGoMZ+q2C47cOjYIKRFUCeKMVZu0LyIzHm
VQxeKNVJMXfaxeyA5irIx0t1HuhnhF35Tgnh/qZb+wmaeJ3M93qO6pIWW6et+yV6O5LVRFlKY15S
P168XpUjfW0qc8sxIwTo0sMcY6qDMkNY1y8RLA62uKH9LgI3uyRGZHP9WZXRK1gssZ1YIHPzN29O
SpFhW1VLV1S6CN7NUOnBkeg6phzAhlkneBUcRaAExHEc1OK4diZHZNXER+2zgNS8ICOTSde21ZA5
3gXSWRWQ6zrUI5Q7JmggfkBknwatmjju/ZMsoiHoV8CKLgox/SensEPu0oOnokzuw7+AUALl1Fcy
xlpTtScFcI7IE1Hdd+jrvRwjm4iwPJPB20syF59m/blgU9zs9mKTavcxO2Z5BGAJbGDRgvmN077L
dkgwij9i7ODfMRR1tHx8G/fR7ocTFQA42cFOpVIbJ1caBYhBJjRuepu9qY6/oQ7xojYFrYZcEQ93
F4F9SjHoXlu01p+Qf8NYSIFoVCowJhRzFvlgOFA10CzhJICQTu/xDLb5wwC3Ha/pvPwFb5iZDdWy
AuZqxIRcCNrBmzXLb7PwHEhOOBxeEnIQmXHzezEBCcDJLXnndahOW4eUUi2lNKlDX11j9YhBvo9j
5NcbUVjqAccLoe15A+a4mMq6DPbkC6hVCzM4eIX0JTKZ6rTMMe6LHj7GZunD8/FUMugHfOskUBTY
vouyCJFb0BRUA5ri596ytlKwDqUEXTz/etLw21HQKCia2FfSyCLcKcQmcMuzA8xnt/mFJ+SUyX4Y
hd+Nmb/NlowiXLcbG1FlpTkjGi7k5vnTprGjqHCUwNOD3WVqyYEJrTPP6aWXUueV9rcxS7+1TGMG
UuBfXpKbZERNwgX72m0t4EnuynCpnxHAeg5DHwfdFOVvLjWoo0tS39IVKpL+jUTwuRSnJcaldXri
xZVDyxa7zk7PM8mklX4bhsRC9Bw6nLgW/Js18MuSvOVAyg8ibHEXErPPFPRLz0p60iE9GOLRZjhO
+Xc4cnnRx1eOIwfGo1SlD2niGDXxXNJSqq2/0WngTc16+SM0lwC6X0P1HsoKbH6kbqKXGTrQ2GST
AEAGQhgwClOWn9PZpLV79YnxWW8XRqhIXNIteK+XQCj447hQAE3bgUPIChv2eQUXRUEEsyA5UHO/
M3FWDsPN0i4MdS6Z0TLP792oHBYOzUctwP/VLsqp7XAnZIBbeVPwLqDyTg6HQd832VQL0ui6yydF
+uli+n3Dp9pwHYDNLr1spoVfQLQzIlOXQal+nXoGCcnuXAtolhM0U0WxhNqsMYEhgMWVeB8GIAEN
MjbWI5MBoamJMcLiau3oqdYIpfv7cNrIe8dSYAHh2bTYoZv8spas5oNbcl5kjqQsrzii0fG7ehuP
8rvhcFqjz1czBRoGlpmKCbAOs9zccHBnUMWYgLUUvSh3OCFUK/F9sE/fDd8ku6jDLFv2DuFVSfna
kaWHgXLgcTi5vpdMmfZeMgkraf1PUElScpbaW8ui/r4Q5PUf76WI+y9Ih/alZANCm06W9pl6FS/6
p0D4G6GkEkg9f+cLW2BqU2k5iqROaJe8Bb5ybsODs0oJH/lEeSV0gpC2V+SkzDw6d0ITf9N4toke
4unolq5FMiac45EtsBiAbl9qdBKp+NM/5v5wD1Kq4JC5BW6rHDMcwL6Wi7G6vgJcPxdtEaeH7H79
NPiOH2YKa3k2uUxxmtbpaYTth1HBRTw7xCTIPdvs4M1TuGS0RhxNHtRbZxf4LtbqCKohM+gSDxTc
IUSc2+yQsB1mh8xGJIxyXjW5Uy1buhJJS03O2xMHdScWqs02zR16vZcVpAf7l0LV6QrxLfBTc2Zc
Wzm23Bt2ELxCSf+1NHFndH6owhHVnkfuS7jjWA5wxh9IjYFqCGsaajdGOH7kHDRAs1XZ2H2jcZd5
6KIbsU2Z/qNPVRVkAeDxLvPb9RS+r5GsWw/smTFXdLn77aw4oUt7NhIl4r8zzx7dhnPLWPwP+2Uz
AKA/p9XoxLJTqonLczsQ3NVhQsexw6FTp1VOA3riVB9eZ8XS9acNT7NC8Cx0+YAxvrEKg2KrqJY8
jECurrIczBiWVo3lbgGkj22gUU7RCkTeHS/bpZ64UfFkTLsh5J5EMj9NfqSJHvXcFfNYS3s4i1nS
34bLpreXWq8Yr7OTjbqTgFqbJ0jj+tFzedEWeRBGx7IA6247+ifnGRGxkYIepF9+WCDKADSD8vHv
mvHKWlEiDoV5VHMXAoOwPbYrO+GFJymM3mkHkH25mTc6NItBnsn5A11Y0OeQ2jtjuCW1ypUQWC7M
hGdyAL7j7yLqp06IahpefUbwzIBs6uVQcX5qAOUjJ7bzAEy1xo5ZUfn6V0Lw5DECsQjosNBCarJA
LPZAplSqLxJ12C/At0MGQAg7FTFrpjrTh/D+GivWL7fjK4TDjW8KF78MW2Agon66Ufy7Fp7m1ZEf
5lBX8BH+Ac7MlGlV93iICNjFeJHKeJA0kewuLyp0g6ZAYNCWaxsIIU2eDO02fN2fcBtWBCaGrScV
6q4RYTH7fJ8cox+QsvQQLQdrexOxSxzO70TePwg+W/KcZg61IVsWn94a8+9V/8YxbFue2nrVRgby
2IoBtBbe9QKoDFH4FSJDQntwazzDEP4GSj09m6FsIdAzRU2Ly4IvTPHUAlo0x5Hs/MKALLpgaP+u
TLtMaPrIXw9b1V/vD8oz+39GdaUZNhcRe2ODqTFCNVkkcRMiY1YLhfI+gHQ/Unpx8ITZkmRlGtrF
dqQwFF36OujQD6VguzBbRc0SV9xdyfUCClXX4pp6cBPHTre2K2hXi5PzDxdQCex1PL6vU+GBexpe
o/aQR6mWwc2tKOCrW0bFfRsQLc75lBeTtF6Zrsz3xIhb65jr+qCOIJrjsAZ1psitoFDqVvG8BNkO
NXCAxNMKoMHiEw6xuZEO3RPf93imauifqZMYYZa97SVhu0UyT5syZNTLI0/qHqm35dPrJj6GJG0r
tArXwDYHJTZDVBmtKcZx5JfhGHDzotl3YUtpZuCIXng8+63epGesEgt+oL2hgkaMxq9JNb7DSDHK
35EQsDl2xjs2njQVhGhQeUOPKXmmBxrOYjdH9DjuSE2ZcnFXvtGVMF6WSkl2lezI9mBaeAQhFnBF
bxEYLq1hIFr8p7/x8Tyj7xWWZipJ+uTnYDTPGWzr7Kf2vb1CEbj620V4yFM3iJedo4YYvMlwdI2C
/dr0N3ir1mAKfskoUFwQDiQgENFxoQ5A7IPiILNy4wg/IPulOQdcisvfFZIQMxBCVrNC8QWmSCiH
K5OTPUQ80sfypsfby8urhSC1diax8wr/DnGayp6UWt+P9BxhtYCkv7fTYglaNEyeiKuK/SrZ+9Zn
lfmitHF+lXxcVbcc560Wg6Ot3YY58Yl4CP8dNUqSQeLcp6dMqDsT5wBGXE4IU1Hi0H681XPo0g1A
vxDcNqrjVOSEXmZCuk1XoERxvcczVxcgHGXHlkmPicuiFKg4ODP2+apypEa647sW6BDRJ1v5rIwD
4nLr0bBCxw/6C98OwYLTTUPKWkQioGQcz+vr8I6Y+EbaaqKI/VGA2gtf2n/wHmQpJTDU5v1Y5sdg
s65MrZwSYsx4ymvZLG966wfvU/uUcpTOSvA1rq1KVNU78vG48t+bqMs96ET/i1G/4Ir2kegw+FKU
dtnG09uakCIR3UJFG4c7I7+kWIKG/rdt1kCOEOzx8uF8A8kMn7H/mTNgKLRnIXV1pncz88sQ8svy
VZfbiPHy9r5DBJglYyl0g3PmjKN0836lcF6YyjBbshlyXIOFAthwA5KbHNOK/2sB5TmYSViMuxwj
4OmPdOZsoHc3aMsIvkSb/zEHJ9reJfgjqrip/BK1qL9okQ8jZo/t+NvsMDcx3vnAuCewXtRe4tfu
d5pBJVPBm+vVUmHC/48LzMNETEGtjOxMwSoiun714m7I5JJ4e9xfb19KVZoFNqfpYBG8HNR0h2Yl
MsWst9gxPJ4f4i98lzn+FPDyXoNVysg6RnNHNwybhSvyYMMO9rQ+bbqv3Thkf19NKFR+g0SyX6s0
D15TnozxowtUtoZQ4HFe5knm92Ha5+XBMbWG7Cy6qQyBR0t/TVzSD1CHXMSYdp7zGiUk1j6VGPBl
ISe5rhmkq6Ddwp6NLUt2GJ2UEa8slGdzRGIU6cxy2UQtYV1pHMJm3oGPwo6Tq30Y6r+TVni8dT5i
2RAaqKy+YYXCxm1QyVdRjErP9fxo45ryfAwugA+DoOQ+hH9xEixFlGGohTEgHtL6rhvz0Dzfqhe8
KrCK5zN205jpmrPE4Uud8JVfll4epvzAdPB2HHWReVpx0+T4CYaf+G/4LSAIXbpu1rzrU5siSbfF
jXvvGxGuiQKxtjLB404UT8k7RgoZt/kvfYHWV95l0aSdQ5xnueB7o46vJV+BCZ71xPYas2XHhnRG
uEv/2Bj3FpXwilZHq+UruIxc2NTzMxQp+eu22+1bleDa59HSyuz6s9hvUWLTvhUIqEKSSqy8obfS
Cxt2rFDE86FSVrAPoaMDTsx9YL26o2mr4jFyUlfuU70iVasTECrbqPKjRDA7iVqp4r6pbjM9JLPB
BZ2Q20gt2OV7DPWyhOM3WVz3fd5dF9yiUSlSzoIOPQXJ1kKpINxLVFF9FdAquYGgtVtnJrNz8bbT
OygM8AcReQBuGjN4AGTPLYjRnvB2j+8fkEpai25HglabDApna5cxrpRcjv4hSn0vS2B12Hh4QmdE
khARqsvMWiPgghcG2RNOe0s6hos0QiY8XWKOgAMGT98rvZt9AvEbwJTj5/qM+1pAESE4X2opBNIo
EGK5RLiOzXQnbhKhwzgFHuvNVnWg+nQ9HehI/Ent7JMUD/fy2q10VP/hWPIa/Lly88+Xw5gnQQw6
U+QT4/A1aEqDpxnN0Em5GN7Gf5hfpjXBLeuRkCLq+kyhZtepWO4hH0GDc7lTyY6NQjAnFmOoCrPe
N2+aHcsq9eCS2KD3PGVcTYXnktcNuHwMJp297cGpYAVMyS+v25FpIbF9KfcVTRcvZmX4Gs0GFkjb
246MU/mZaErLArr476rStiw4men5oXCduYK50nvRzd7GV3+CMucTXHt6Xe7f+jgKfrrln1Gacewq
JbjLuqlUVgmXOQrRtInFLIeGJ55C0ZLHPPII/dBrOaqh3c/S3eWYNXN7S9GKNFAVy85P/g6oZGx2
QtovLLenLUQDD9SPr41IDtY/Aen2N8b21jfW/oYhiT8rORrSLXz2h5EVFwkQIdy/v1mfdzHH+41+
GfZkXo/n8aps1E4Z72MAvK/7Wpigv+K8T/Gf81ppNQnixL4TUEUvVQzABc1CMkwykzxTpYiz7HDp
X30o2W/vfUw9FWAlwoe3+F6/PmxjthtvOTrDyaoCtxDjqJcOvxVJz3NM8lRxqpAD1iZ3blBPxaZh
2x6iEH5Q4aO6BOTzOQddQYBTCDcu9pw1leZg3IBWuNExBwNT+EssTITLK0Oz4VSx51qGBx20/CyI
y3gomiu7vVxw/Q2Ghd8eKLRCadr1RL9bNTpe4H2OFm7NwVyju/8iZSVXHyeEyOit673AW7WcE6HD
kulLRBEoGWYb3ROC9F4jE1cnCAYVQYCQe7hVCVZw7BtPPDUuIBcEROre71dJxKTCbEMk8son3ctu
NTeSXKpfyLWJl0l+pIiPiGw6VwlhzO2QDvwoSWdoxv2uaYj1L0d+CQMmNpdIqC7MLQh/KHoBlrRJ
OAXrYOqSrN3OQRDWx3bE//aRluAQxVsTtCnwv+/8Pvd4J0AV/0ClLkRKQtLNDHQcvXy4cS/+2Vh0
1Vj7Sb/NhirAzRvguHTCyHbkFoARF3My0zIW2sISt2i4r82fql9+5Y9eNDMOHiyRVB0Rsk11TzkL
gA1UIbX1vzLZN9tFM4rcmaxwgGn5VMbgjJ/28Xp+Uh5rWqBcKWNuIrjVSCE3TYlb0C8PBMaO2FsI
J1+VQajf1oTq4Oiz35vnVKAueiybOCbSEjIy66xmUgOaGKrt8yS9dXO/6olKu1vQnHks1uJ2QW0X
J5Kaoz3XjNtFE/XAiiW5W5eIyp/I9RIpYIAaRRoFGm3Ct1ejztHdwloelhSUJ1200zS7mXIEkJ3O
bEraz5/WZ8QfXPwOystHM3HI8wxTk21FCH5ZW5E2bCa/RmkdwSkrKNHTie2hAuG5vQcjUAGAUSkU
A7rUfnjk2tUa8vc98n1voPb1R8YKOl1nkYs31zZfh6eN4DI0IcbQHL881G+E2ji6YErkMDD/UBeK
u8jfxAdF3ubE6xWPdghvUNlL7ZHE9m0rAv2HzRVq52jD6/bQ9ubyTpLASuzIX7RWjxFEMPLo2N45
k8jjPgrx8JV1VEBahX2Jd3ngvaoBtdde6Uz+NkCw3HVAdi7bU1TPWLcVZSLEJft1xYf/fRz4AXns
lp/N5oGHGaVhVjORvnOivcN16ZU/NwgJmukajtjyOV2FnnPSMUC3ZI5bcvviB16cAeLsv2y4+be9
1UkSChtGAJKumqgJoAOkjXUAiI+9EDe6PSChb8jAxXp+UMgMG3q/45scMwsfBOfAW7f3zhtaijm6
HB/mPffGFJeQ1z3cPH1QpcPsHA6WqenU7Bug/UHtyUNmHVzHCMPnEZmSPBnpi+uRdJrlAOWYQkQP
BAYjJ2KWUXWq5Zi8osT0WR1Ea3mfrLJ/mcKs3ohhbNnH2XmnT5qQCyaJebeohX3NdYHPrWQS+3Wa
Nx3PkmysOAFRf/9iX1srcpkcP94PgcrSE+hgPJprrx83NTm+yUju0OtlVmeQWIS/6Vb7Yh6nG1s5
xNCnTiv6NuA8Ju9ZqZoF7S2LzHyN+aDwiBwAya8JToKyE8HU0fHcSg8wbSl72FYd/PiMsSxkJAs9
KShv/C7wQoNchyDhDlGSRbAT2TRufcm751PSxJsoqHo22bVOzmLQw+MqFyur8VmY0hu2F/vtonGI
Cz8le6EyVwsetdVwndS49UsQDYHI4Pa2BdX6SknPa0o+SnO42HHcyacOU8BgHyIMtodapGTOUkL1
bZAEhxentJ0/3Lj1MubbNoi4cPvTtHjVO7AtNP6xc3TMMbmb41OnI0pgBovHGO7oZNVXuF+8AFWh
tGZKce6zUZyqj16yk5MQ37sRy8+tWRYZJbgpl0nlgeyGTsw9ggQyTflrGvSsINP38SzNZR/Lqom4
dgaf+wFo2ElxcHCouFPhlRhEiUuCChua4/bJ5Hx9AGj7huRBc09VS2haa3mPXj631O+uU9LK6HZZ
pWNkFnXLbqFpduU/JQUmTYR21SNE9zgMa5z13MM3yO9nZmbxtamw91Fnwr0HS6PlE65IJ8ASmXXx
a0NmSaXOJiwveqm2D8vQrLQ6RolvWxOaKqlMZKRtSuLaynHjbbzELWfvrwQJA+B0po3l6ExCdk6w
KzJ4q3Rk41UxrZl4F88PFanAeS11YU9xhOB7YTtQ5+FhFT6oFYdma1JrZ1v/q+0ctp9U+DeguJuY
vF4tzEEiK8jId7FGTf1qib148YgdfmWZ1qAjyFpuk1Pbj0ojw4JxaDJMMehPrOIu3p2wndk7DYOU
lp5jVJ20UvHRIDlyR31ffuGjDZvYzUYXA71BSGWAmxBHMc2pSzh0CSZQwUxPl3BHspclseqCmeil
ceAAJF6QLNEAAUvaRiknVXskx+hxciGtfF4X/LnoGt/7/DP6YdUcrvIISpH0aVVkXVcy+z0R5l7E
8QSn28531eOI2gHKX7wWraxwwQbw9TFGltX8fbZJ/jWuA7wjNEGVJZIDtDQY40TR1qwjvljnIm9T
Bp4XMGWhcCYULI+AEz1ZpaMnFG53j6DQG+PiuoMjKwq5ugLCRFgAwmZq4PSkRUiZO/70ukckyZoM
j0aBeaFIi6KgGMz2uICCAjXdzoB+v0QH51jKJKwcjkkjEbv6WWSxBHQFGUY7GtEIz3yKZ24AokLX
eIJFxJPAUVv3iZvovY/MjHma7gcFl+J9DvkzZUkfHUq/v9+S0PS7wXB/wMO77IrQ2nrK3SnGmv0G
8G4bLAxFEXOH9wdVOfKQr6eYFrbWGr8bSD1PrJaPKhwAEvWyS5AOn/zVGr51/3JnHUzqdmS5JBPn
p9AuA/eHy1ca2AxR00KIIICAqmZlnRUK7Ld3iNpYTLaVMP5KhLMXfKWCZSiYfRNzt93BT6n+5RF2
1DzJrbuMGgJOqkYJPUPFsOr5k7zl6tVV5QNtwECSLDeYz7msr/AcJdmUevM3HbDguZSFkhpDM5CV
Dax18ZNi5oY3v6iawr7KxuucopTyZ+sRLQVoA4l2pjLoTY8Xl3OD/wyRlS28nd2Hv8vKT9opa9jJ
wtlcOT5e+yFc/PyvLmVeDACckj4I0R6Bs6eR2SfiXVbUN3Yd0gYBLGOfmmJ8UJOqZ5fd2Oh2rq7U
rgB8ophPcyurNOXlqElgnx11s6zlkJqA4oLnwVUScyE6McEVrg0kw4TSb4CZqtMT4t1/gfl8ak0c
Ap+v/FRGDamA7uHkOUu7uwNQS3w2t6F68XVGVUq14awbFT5Io9QlxLCTOv34/ZmZ22AbLXVW5g9w
yzDPE3jiO0pwlY+g6W/YHdCnPUnF2ldPemejW6LEABg926t0/VlqzDgTd/ZOeK1v+a84rTU/ru9k
IDNH5F5Jv5VF8o1VODZ3/Fs5kMxedSkd1G3Uve+cSJWGseASm4L15gDuMfBKYmAIv5P+TpF6HSs+
OqroxJ2cNzJcjq/jAMpWv3qDM7T2GhmeUxja78rxxCheyn+MRYxseGtaWomUTo+XfTgu/moECMbU
tHMwCMgYRavPs7tz2BVqv+D/kffGC1AMTWAIFl6b/RptV+UJkFuwxmnBSUY5CGNwZLP9jKbn5ekh
135Mln3poy16AF6THb47uEDOx72vM/FSRAy5EDjD+jPyHrLtwGaxgFnHnpC9W2PmL2NSF/tCoGnT
zwCgQQVVyL8sV+YSNgqlsidiXLeXLQemrs4aNsEsCachYL90fZGS0SZZvohuo26IPm7i5Irloa3q
MRSw3yYVsEj/kJ7fAba5lrRZiUE/IzN2qHTJXkZX4bESi+TDoHRw7ZCpTBDhNdM0lYLFN/K0B684
NJ5wtpJyzsj2cFNDsVCLGBZtdVGVAW7C01bIZVcKnmvFbgOONcDuy/pyOwFwtAhSTwnT3X8R9BUL
UR+fEo67N4zDHr1vcbmZH2+bCtVqYBwGt+7h1vNmYfgb1gAgv+mj8JGoIIp9Gr+T/d67Crdc+IB0
SXz0rcx9p2t0/UsSHuP/Go1c3YeYpwZswRJutgMqvBdm1faLvlnwVMAstW8TmQk/WUX5C1osC2Sh
KBRevobhwpeeRun8CdRlQ9ZJ5vPpSmvcKFPRZKtbndewg0RZy1iMC+j3bqsc5Huz5ECcA3eG2OAM
qkBxh5k4ro8auCvfSx1si7Pb3kNffgQPa48V37dXgeo3yBlUk98k8iwiL4xs9BHaBJ1vf471zALI
sfILA+SQNF03JjPdmwc9s+tv5fGLWcIpQhUNGxLQv1Mwff0YoPDdbSJUwp29/GV4Mi9sYmuRx03M
61BPB8VVPMnGlH7uoW98A1EUwmG4PXF8egn1V937GpJ9GoYqSqvnyONP9S9Eq4+/cg0/qeN9vDea
x4ranOI3P6ClZGlh1OuO2gKHb9PYthwn88Kawn+0oXkx5K5elO609YZXGLQVxVLDntuI26p9p17/
3z4oq/Jky3AhJDkTbxmiwbB2hPV/UjUyQga/hK2w0bNGnMsEgh4RtFSm1iDNBgKGrwzQ9K006Mtn
2/vzquorORbGWPJ6s3Z6IZhETlQhQ1EMaUxj3/4isHuqeTFUUE5gbKEcOwB9u9iv5sfNQDImpexd
EWKKYEegilYn9bhFTn0e+jEJld0WcP8wWz4iYs27yh6ThwtM2kIyF5MYG45M99zM/hnQnxSuQcZx
23W0Uu6sulIQa6Uw6pHqkVedls0G7IMGpnFP1ClkE1AFYIVQ3//0uiKl02LMHMJiy8PoDmR4Fufa
6sZSPyAzQN888GFTEhy7SZ1Bb9iOOM60u/Lu8LhLY9fiCluq+H8eCNIl4j50i6J9OS6eiojDAMaU
ndKQaSrwY2sIEERO3FytZOgRD26jfTlY/IvGow/ChZyOO0PQmSrFfBfCz0usyZ0Ry3+QaeppdRhB
i4F7eRSzViJR0RTl91ErGu7x8dkUtMOB050vzPvbdYfibd7blz4Il089j0Pq198PjmxSiKbcr4Uh
Iddf9ilhPZIABiOarcdIzp06bpRudSbpYYQxf9ZwZ0sNRNQifpiZ1DrMQ9w+vhzOpNfYOSTWiqIK
K+O+LSAqz8g63U1RMdHiLhy6N68sEJuwJ7ZfR9a9U8RPPiWkZNfQR2snUs0dBb1GS+zZ4yeQqp5p
cfrzr/vCzV8jioganXY8L/mO75Gr5QoxVCiKn+ToKMOlokpuarTdhCA1ppPbGL3Crjm2fkCcBLWH
+fWzix79duEyh/cQTtnU+mcwpbpYRdyXHwmhkovBB5B8A2A5z3fWHROFC0LbHa9ISovbOxOeW5Ie
Ap8EjvrQQayvHkLIO7uPlaIncK5IXsyHpY8HmnzSDX1iQPbIlXIdYtumc8elwqZJU9o/HhUAwZaA
tCSRcg74V3vUhyjnqDGO+v2uJd66OkqaKv9M/P+ZGdEItgHA/qYVYtp6POfMuA0Si4TREiiCfjlp
6VffFvxMhwf571CpM1+8MEujTIk3a8wAh13WSNdOuYVp4D938q/v1ay6rA/jE4qk1ThewqF2sTCR
XTnLauxNRGiB0ohE/mutpYx74VLsYKv8XVTkEt+MS/bEKXWt5LboexOgrpDbZ2rYz+mwVJu/2Ksq
9QwdxTtJkjN1itYmDkdorT1EXmkL6hiUzPviLmkkkGsOGGuMyM93zoeB2X7vARpCoDDGeqVbRjl3
vAuopUZU0mhlFsv/2tPHGiycz0rYqFn1yFe2P75xei7z/MpwRryCSDcl4CJ0FV7ffgWTq1zA/kQc
1M62N/5E8UD0kDxNaEnT5Bb27jNLkeqfW47ZVThazfVURxo2NCPZWoBFDuhlNyLlp/VWS/kHPCWK
7vr7W7FJ1AyisvRCdpKSc6u3L9TVoD8bJSg1NxoNYXal/KA3qojrKT30ZAEQ4iYIgOnsfE8o4S4o
KWu+t1oHesFxdjy6GLO3O2Ht1epAys0l7HhvXsdvRSurrTBYNSDmT2e1MExPBodnySX8Fa/2rrka
saCxp51NTYsruqt1rR6wLhbgP2vK0lTffgvWw9t3YIHkiSVQY4DvUON4xE1yTi8OfItlN29di+f8
1YP9i3FzlPbP5YkKGhjqFDZ0J95o29+98TR1dihbKnMqN/eJMj1zoBPMAr38iwBk+XQ1Mxqj0Jdr
O5tlvbPT5p7lZhiYJZBn1u1uV7Amc+gDNWUPb+BJs023lP6N4VfyUQgM66odC7+S9f7CFdSR+s5Y
e4NPlxbotLf7nygP2ixExj64xeuC0RcCuuFgWd7NFkjhfkKRqO5k1nDwtuJFxfyZmxhJA0qBTjrj
WhcizOFD0+KVNQMJKD20HPcPKqxWieIjdIkXqG0mxndXRW0jJtBTiElGupUhABcV7Qm+9yymbSpK
tfGiQy8X646tb9LOoWAkFk7sdtubYKYQ3gpoU+TEXq4coxaMIND6z7HX3t2wgv48tmx+P17qpzHw
fI4fQyYsfP17nhS3TXDTs/eKHWAH5e/ej+P+LsF/yC2lQHt6BsoCCCRdfEgsKc30GDbqt87KtwQ0
WbChYyiQ6FS8ITrmfLg3jKyeVd56DbwB7m/kRUJkttifLDLAO4TviiEGG77YZgT6gqQ+OO/0GXNz
6Rr9ehFbxOvzS3w2rl9KuepqLV798IeXy5SUr6MV1H9E6FnhtUKINtp2K/hwQbW/IdjBdryImNQd
HRyGMf2nJB3Qjb0e/KqEsGRPgaSy4B/3z6UwDrrlum2qcByqqJrRFY9EuCrYaDnE3x+ytwj1fQQw
azgdMeSdGkFmQo1CIVV0QaEQ1tZcRL174cZVjXz49xkPGf3AMzKf76YrLRC4E8AC0a+noWiaS7mJ
xTPLF5uZrCHv3eo5rLTIVEaT7BqKFKbLTFd6yLO1F/SvpNLDoQGKMqLDriSJ3KGbOcFoxf3yIHox
pJBrYjj2hX4Aw+PqHzM7Sz2Pj0RAcSTx85Ia2qduljZJvpqhnXzV1Lu/vmlMP5esOAusMD1s8+bq
x61nRbwqSavUI4DYFWn3Y8xqP9J7zgnEyRGlRmRY4OxXA1yRBYtZ0VT+8aTnnMlUS2G7J1ZYsT0b
emHrduE7gk1J9WMV/17wxHQTKc9OedwPSa+/EbJ5mXGWOuMS2kyXdtiGVtla+diYN2FMfaYjrBSs
P3WnrHhrVsuI9CAV2TWtOA8x5OvTGnbv/7SYA0/xTgNwWzW36tcpYWhEXY5LDwWusqQ3suV297U5
qYGWm0dQvNKxWvYkSCfH4D2qZpJhMGY1uYk1p+/hltHDgE1Th1wljAAdntk5ZXqc5Kbto99Ogo/s
7bL6IxIgOlS2uGqosylvINSoSImcYzQkESdV9eukZUxmzqJimKLdy+58xdlfKpe4rHwIQFCxPaZQ
EMgihFINjstRLP6rABOpa/F3cCTXsR5wq+PjiKsMGe+bBumrsmJ/dCtoiwuKkazySfdceF0U9819
ty/n2dsBSL5Wl/CT0+Ekojnk1x75M8woXxF12mPh4MTzBhghb240S9MT1jdNtnI6m9DgD7lTUd2/
rWSG9vTBqEjUj+r5EXAOdKdrNeRMO6X2L3Q20PJ4Kp3w6tYxvB/ln1gh/e179d+2g6T3v0W4EPNq
DVZPJ1rY9GnYcNmAXUBQdlK3hhSkk0rpNYs4cXVLlrkjTgOLPe9Y3/MBd9YbDSR+mL5272oRsBOZ
DBIysHEpwwCLLWDssZXeJLfpDTwKsqzS5NvVYm9wRVUShemWtqmy6ZcPmS+JW/qEMvVCsP2GhUxE
PiGNPThEcxH+OTER2C/IcUWAG5s+PEm2gelV1+CGVZZK2W7sQipCkz5sZyRNWyMCX3Gtz5T9MynW
WbLA5BLo8cPZeXR62GjTrv8ei19FZ2bG8ReG9MC4e9+iMJ/d04dIpyzPoulwt3FD+yz+qOSCBEsq
kyrOm2stpia1XYT8KXf+gIDwwkIGoeuLFnWdB3QzLBaugiUxn9Mas4tL/PZYACfprPE+LAEtXbeL
s8Bre0D3vgnoVSJf3m2qbVjjd092gK3WAF+/O4SN78z7cEE8vDvaax/aHoRqGVVZD8GwMGa9JPR8
ncWmeSguyDIDowwacUelic50xWlub8Lxa5yLfLYHYwIsWWlWq55F03x3osQt8XSQqGQNKPJH08s8
y2OuIkCulSpEMJTMJilFmjx5GmkTeWtY1SkM3Gg/IWVsvbOAys80CowOF1Gr5mC348+PEZIWftwd
sE/6LU5wjvZYce2BWvd6+EUobzCQYLEsr1A/I83O4f5DaLBaNJtM9ffXj6Zp3HC2LDHngv8rU0WB
xlTGpkq49z5dBH/PpEJb6BvQEJ0OO7lgtDkIa+sHdRd0DBzgmNqaP84DsqsdEug2rMMCY7rcwAHQ
f6NcfM1flC3/AfV4vLh3iPH04XomEumX+Fnx219LwiCNX5unzj6lw+KJSnSB0IRpym4lRWI2+s13
v7bzTmX4bKB7ZgGV3AXqQyW5rezbKMMMFBIjdSRpNlF3hVhGCaBOAOvTJkzhZiVENhUzQVWYUm6Q
0mmS7WRyyaKhKhHWs6/oVG09tAOlbVvCePRujYrWVrAn2PRTOV/RD2GfrxsdE/BGycYyKw/OcKdO
8oSjOFXpxEaa8jdNyQydZaroyBw8Z/7RHYY3PXWz7HE/EV908U5hMi4NG4WaaK7EzafwzZdP0LVV
SPr0ACUaFVuznTuzGNogiHShoCnwDp3uWD3Eus58pcbKJ/lZfD+lE+9i7Ay35NdlXdBZQTTszsZp
37u7TWVs8YEGFBJlXGmLlY9+sMMax4QVj94SLHtITd6Vw4bWUJf0L+7veGmAtUOmI7V73QFwTE76
KCx0c3XAhR07nrao19MH31KDTwzoOmH9MlPf0tVig0Q4YWUSK434oBiNOF2YUgd4/NKhIP3A243W
7vMgmYO9W6Fz07SS8hjVhDyY3hN12Z2LCL6XWcTXYGAjiVpr3h7hu7K8CzSSIk5EdUNkFCN/d8rx
9JXhJGb+qGcvP3+YW7trqHhe3L/tLNUJ/UWPIj6hi2bTcxDSAW5X0S+9I3H9qOLcd89AgqXeaZ8b
48FKFPwf5xC4+v1hj3Ur2i0A9KEq52EFEornLOH9RPUFjizKYTUHMgAFj1iNyFMbzxZ2nRNZbNqa
Dqtjamq+dkGo0n+m/2rVhaccQ1MQAC4pv5P1Cn1xP+AFpuJZf3YFakUoHcmGS94+arMIE5DhNCZL
YpWyIfII40JwSD5LcjU7bJ3XNJkESeeDCWI8HGxn9UosI3uxZDbEpGTST1UOFhPRb7SQbdUZoJ7c
o3xkSoOTbXVASt4iTVJiIISJIyWSVx6huJ5hBo3dx3oJDWEDb16pdRUe+DdpDcKRk5ZPhDegLQot
QSEyB3vTvGlUF9T+dkWVDCJvD8W6BpODLegC5pNersaztAjmT+viRunMdYqCk5E9YVZzRe5fh4o1
+XSiNP55WEM9qyaksmaAWlxw7IgOjtPfyBTyITNK2NQ/GhmVKpfomNIMzSfN+uuP4+PNspAUmZVX
SqjfGaRO9AvFSwHLVCIlxRw8sh4RMklZhYedLwLA1tOXP5/ff1ZUorRNcBfsW3B8VQTqKXyNkH8d
5QKW0Tv/65NrnMag8HXKnGTGxBdk2urfEJFPI2ok9ejT9g2MbmLqfFEx9p3thUcaPT19wiZ11nCd
UnAvJud4Z68eTJHgHaXUv2tlos/NP3AOKVlMwvXQhYxvcrzaaDR3hzTR0sJiukP8DcZ9yg4OET7U
+74Q0d8XenOKvcmxZCqWcNgCPNjNpBQVnRflp9Yin0L41eWCbrZ7kRGbys4B7Blskbp1vi272fre
W0FjBsCTKeOwHqf4pvqzn4xNFFF4XFBhRw0DcNmeUHLXRS25FiqjEJinucmkBw2Stzb0spZrK2ul
E9ZGPaGsseh3EP+YZmWp77646+uPiEK++DVTedYTuV5oqPve6x5903DeUah/vofGDS+Blip/nkCP
+fFeF4CuMh6h4ZIEhK66os1XF6vz7EtPJs4aQOUjIBIOrJ/1eJwTBmTCl4prEjPf+uEpHiMgjalp
9/DNBQ5Jr+hou1UVjEq/OUATmnnIQXJwyJZg4tAr6TGhvyr/3f9IeJv8UQNIYLAzEUvPU3rTmV4a
ouD+po+1HNa9hsX2DPjHEoFRZe2nfeNjsWK8hWbo4Cdo2jXEo6QhdCd3ZNaygoXtX4ufV5CeQaoB
WhdwCt2IG06ZAMRzupJSWosRKzUX+yLzuYvMFHVVv0MhMi0ZnFmy+63Yi8sNnZ8yrpH9/1WukKmj
K3HEqEk9WjNhyaKrTNuqu2UqHvGlGWYMWTnLh+0M5+RMIgu925DL3kRkLeDNBn83dnujUWLf0anU
vGCJmPCK395XjqsNTWKE/j6YUaI+bD3kS1xelR7SkV/vNQy3mSkdhQ3lDAOWiJxI5QX8HlMaeSvG
GrzYDj0NY64L9ulSULg/CdQz36hMnmRlUkNv6d+qcwQyLJ2QJhTcApY35lAGCDQ93IFBeo95XvQY
/OSObMXSxaatXwI5z8kWee+/bidB2ozJDaaxLBkygRfuuFgZKHg8C0bKLzlBBXDURFQS2eZV7yri
1pgAe0sLZI1pb1T3CQH8CPCzlxJfbQ4NtunKr8f/U9k1kbAEQX+gwmWwj8numsZaNGHgAArH6oyu
2ZAf0YNH/4KexOBt4zO/Jis1m5+V27sUkHnw3T0w0Abhw74OT3sVeFWEj6iAAknOKCsmwRqqLGoO
PYF6RMpqvNrgWxAL/se9GvXUmr9p2xI8S+NWguzjOLWSaxZHchQOpiuJvngXaOYD6ieYfCeiDB/m
XsajhCYNFpvN7LXWXY5r4hARHAVeSJeDD7NbTUcl9+66/9Fu/71JbWIpCOug7nQ+e7ykFKelT+MI
LcoHTeCV/sQqTlj3AUduiILsB7eY/0L+QAk3kupZmprgPc5pSzI4fKs6AQTxHHfaVnGG568KOMBq
8ppQJyeznB7KkX0nvIehy3SAJ5AkrM1/2XxnwUpCwNYKyATDzWq2E2fFPj5YYI/38XlvD6zqmlJj
NOIBx5NSRz8OmA4HdX8lRX8O9pUmlQZlzHJ8t7Sk27EsKsvYHZsjCwvWEmZ4QWJydu+Rb+RgoXxz
/afurcdm3cUnJF1b6hIqywxBDZvp55wekKOCbpxX8ngP7ol6t11n5+vDwkcKHahaj5LtrRxmC2MD
nq0bSxVSmChE2TrDhXEbm+fYOJmO18tAIVVl4I2+41AT6of9cW30/srFy8UihZt83BIBTbLpT5bq
H/KTuHuFZagjz2NPkPCvp4Y54zWfcutvsqN6qL+wFme8bysIJLL2+vRB2vE4E+S3tETF5Q7UNrmI
eUwGRscdPwsazDg4n4banJi6RA/drXH4PCp3/7tgAnRVeg56hQzTmb1/47Ohkch8JCQXKsz7GL/Z
OWgUHPrJtVnSzaHAc0q56vXHC0ykbb+BsXbVzIP9ceazdMRNPuh4heNwJivUp2WF0bKLJ9Ilqsgy
QKoDNuSEVMrBSBuXx1JiDKT+VlUTPqU3S9REXQ+fJ4dpNdlpcsV3fVUl8NU0hpncnEjjPeVQNurR
e3e7Jyg5d9oigzi90jtVtjcm841RHwdtfEvn9/zTlrupKxRpeZfGqiTokL6CKVH7ehmRem1bXI9K
5nuNnR05d1/RHumpYJDq/bfXDeJByPbMkvtpBnwGQ//A65mr4nhlZnCXT18kuB+PSeDmxPxMO7rV
p8yZki0gVOlo/5Nf6hGjLNhtX1tBl287KBkAE9vJJwPaM83XyYWwiQLL/ZI4zLJ3hp2PkiAbdGtu
dfwKMElvqiKVmS1Bj0ZqbPbIMxUaifd22MSGFl+JtqqH7UwPpNY8h6OLRKjmZo95H9oEqkLMbSI6
vfEsFhErctTDMrE4ROHPNb9hjANei1jKLRkX/8n220BrQSUQB+Sa4aJRqo26cgkMHtAcxRc3H7Au
7BvjuApqC/THHJkYn7m8PXJ1701ihCHDZMmaAbdcWk0/qKqn2V4YexT6qvC4+ohzNg5pCAseOg2M
RJVywi/9n6N2nsyK+ipBQ7m9Bkj6Ywt4QG3IieQTR0gA8vBiE+JHeVn0MhQVR7VwCmwtPnGRxDtP
pNTl/0adGIyPWNTD7w+Bxy5SHpb2KiwXbyPGYtQLRA7oKIVgChpDc3CA6ArLj2aLdZYdL2hfAwJr
Nm+r5brXs49iwSxC7Mssj5XreeSsHYnV+nUT5GjO81S44JkzvhsgdH8pUZh7QnAXqoRY7OV4xPwo
76fAELEGlI52YOVzYw5xdIZFFIyP4MLvpmF4b8oAZ6qDpWzHBLJEwznQ2gjXrbiTBTn4RQtOpIHg
qN8u/AHaSKEFs0YTDVaVDp4T/b1JJXvFVrNRVRw+bE+/qPyHochf/eLPcwH9rHUt7ex42PvTmn2r
QB7wRMEBHbbOsyr6ZvTUJPpDZsFHWT+Y5dIK811IMArtbZiq5io82TrpWtBupo31lIJkxhIKc2cP
YaHmB7EEiesoKFGsChJz7d0HIe42+Vmq7S8x1MkYadozlPwrFDL7uTdNzULw5gyIvIijA/bj7xZF
5Mi9ZQhgIYhGBzihRl0FI4sEW0Sg0vUJM1f6W3l3BJ2/JuaMvBOcYaT4nXQul2KAmI7GlHZrP6ju
eel83oMTojYVdK79dZggixF6rMgFOaOzuCk9kKnmvdVZRAzFTUjvjNgnYsbjeyEdJnLVbkHU9HqJ
1F8MEXZm4+Y9SOYC1ExFbqcXfCo6vzaumN94IhdU6G1NuRXMglg8oFQjU6NmYgHDmCjFwhOVNx3C
MEN+osGOfgDVBQRVKJ8oFi7Y1tSrxd/nr9ki5cYXQ9aNAMOtN3RWaUMK6Vwar+7QfkQ4e5rPUMP2
Wa+G+DbjuO9b9ZZCmxbY7JmVyOyFq0fQRYCQnbL6P0+BHAdNlDH8ZpQJ0o+EjBa6/7FS68PbwnIk
UprampmkTk4AwOeFbDhaFEdqq0f3j50VCBmNcBS8XyWctxzl4uiSn8tLI6AVsqBk7OkCCjo9JjC+
ZtKvBoO+jCilv54inxN+rW3DX9nxIvYjY/2ClUDOBvosd3tpEy6L/yP/Yxkzqeznzw0i1I+tiuxK
x9Tui/HDTxLEUfDdpoEISntWMBIpNC09eA4G4UuhzIA6R2d8HtG4FhPqKKvAcG6pUW4HTTtxR/yB
sq6sTA7pd0JrH/5i/8GQSaM+NCGYPz9lGGGpK7+Rqz6+kiOtS4XlVpsn3b5MtcMbMM4YcHwgRnwW
YLx87qzMJp2LNSjy1Cvuap1VG9wq1XEjfcftnRWM8jIHOavCV3MkpjDudliS53+4ERql9nNlvhb+
GGwK6csMvdz8f/d/NdpIUJSSXrMXGfR/GpbIfCsZxGatWrz9ZCCf8FRMQru9qNRTAudX8lycKx+C
T5dS0WJ8irl5hzX0zk/rSv1TItEXbc6uZmxxhRdiJfiQqVQuz5ugDsaPBev1jD3T7qaYbaxZbfyP
3W9CoqOg7gwyb+cp9+CTEQxZckc30Qd6PZ6Azhz7UEldC5TgbPzLSTz5emoAybvh9bZSvtrm99g6
hf0nnkb58CDnxMC3dUOexxcGUTfBNdUUgOQsyDxx5RdiruDsKsymVWTPp7FeRRJ2dgUk1lp1GAnF
21kpJx+mYGs69e7jtPrurfnU1QCwjribzHV0Bzn8vuoRQ1uo0sh3b16yggLV8+JGQhrcIdrs3tWM
1BCq9h6uYiEf4A4KTiK1pSvtLgcukRmnCZm+JvzfKvSVZ8ePqZ6+MqjUMA8EmMDlmsoxiTtn7DXz
4/MIpe/WxQh4BsbpW+p8zDNFzCiiUOc+rGvgnnvFIyoKNhz3WZhjA0ZiSUohSt94ANFQZk33kigp
C84ZAeJwkFfoiwaUaJLIf3oK28hKJpORKJ4Yl9NeWpr5lxIMRWNpgiloWZeLrJt9/1XdQI0L8RJn
c0zDf0A6fuRBo0awpxxOWmfzGGJ/zeO4tTnUzQfwOKT1kq/UPfChfLPohwHImBwbC7uv3TOkSs4J
PpR7kcicCaWMoWkg0owlG9h0zQCIbPjtP5Aoczk4jzlNZlv01rbr0aI6u8KSJSOIoUlZV8+dNg5/
I96hAq49gChXLxYRUJUBiKm5Xh7Wp6k7khIuTMS4+BCbfCzTJQ/miQPEBIbxxs22RRVi+HhRNVUF
Mo0upRI6/+5oECvR6DwST1CtQKpdKppE2LqaWSndgFDj9+v6GJyDvTHtmyddNKXS+DzT4fp+CJRG
MUMnV5cfcGiYKPqY65VOOMSV+LDEXvZk0vqQqMx+j+ysw1FKA9RnQcn7clfrZNbFJggtu1tCBXs4
NRXLWJkXeON60sQVyrpTxVwn40THmegTikjet7LI0p2jHU+Qd53GPHnqpMtmAhA3dzG/YvfGMJJr
q39A0AOOx4ZIPEanLqapKZLhIhyywM5vcGrI3IPlwE/kaRRSvh0cS/a//4WRQryvj28lqg73XUuY
A8yaGDMilG426qLT3diz4L47uR5Yq6qwZbAt+QAPTBqqtQheVbj/eyGklRuRCj22IeuhcZBsHcYJ
se/4a0kxEUN6YeqOKjpW831TC/v2NGSGGyDzii1vfjwXDUZqfh7+GBDa9f+jyF88AevK35N8gyh3
JVPzKXLHL7G6RdGOLsVw0O1aOhl48Ez54v1C0jDWxyfmebN4lxLt7dwHaZUlLd7hwvVPCDTTS9Ub
XI55Ef7dxBLnYwMn4PUJrp0K3zZaW3HYHUhqn9BhhwIJhcM+ccKhZXuhg5VaOpzTpIxYAfZESwuE
ujAZzbSf/MEsRMsUvK0kx9BBaPYT+YAqu5FWLHBt3SpXh11fBX/45xCdGGCp8Ie8i0NHCgudJtJ8
ch53+mIrbS0MBPL8uEqdaw/K4BqdctLTBWP0Z7dXX2u9qQHiRj4K2MeLskquR542XqIxfYZrtafy
CHqHyZkYatFu2p1JJNlWtMLAbUj7ylKBwWTyhKA3NTYkxOcocIFKl++AgwN/0HXK1irhN4IyBVAN
mRhgINku2aX5le8XJZWbg+zor7FHqiT7jZBtPp7SQGTqnfchoNXdOM4amfRok70ppTmNe5lCMS18
5G59qSih7PKkUo9e3OwR8Sf6FLyBKbXfwTClvApZpoEwXpD13wbpCwzECaUtGx5Slmvt0YuXzVHj
cvUcRtoWwhPjMrxy+WEnPY2eo4XAuUBiVDNE7W+B3gpUOzdnX8pmpaA2BoxqT/OaE8foHA+Qdh/X
Sqc402AW/iCIH5wStpo6kQUfgN9OkokViVCDO6S6ATItXl3eNT6La/2J2MBQa4xUov2Cl+ly3luv
EyJ90sIuh6iXQSIZ1YMnOsGbdDXU0Uvbs2jqp/3tGFCH9RpYYiVYwTGcHQADnsF07DhGz73iG0/k
2MfYP6xW7pM/Ls/Qze3anZr5PQ/XdIW+R0TYUV/1VYRbIgrVk6ozp1tX3CqSFnENfrFUBvbO6QIc
WENvdWNUO/AairvIoPc5KUUl13lhGKZ1Rc94TqIANagAHqBhyWYAQ5d+q2rMn+UZtp2ksHvt4skw
zlXP5cezdBw3a+ZDs790qM1hLQlsoSKyGcy1dTjPhBtEZfsLIpzYNZV/Q6zR6IL0hy9BOEoZv+oA
LFk/gQg+nJv19AtJaSyQtcm4lT3Sa16jFHOzWKkYuIpjvLvZJiTUEunKu1LIiEu2Rg56HcGGKMJ4
6BhuY4Mh9ziw7N4AmbrVr7SWvdsZb72WXKGZ2wUmO5frBf26AyyPo3t4lnpGbNOY46YSQX5y2lia
ZG8Al/dc1x2pGJLNYs6n2nGsx78MXfBZTqu9gvC1tOr/wHgxFuDE19cx6fqU/ggOLADByjSd/STD
hUTWUKNSInO5n4S9/J8hHs6GZBWcdx6LB8mh7xwbKrxXr/3hrJaZJZPOO/sZ6Hi5yeDHao9DTC0f
4afS4kUkYbkgsQR9cjXTZjkQVpIhKAPDfd1+vaQpy/BjGyi5+zQqUFRA04QMUPIyusABBPS6SEAt
96OfvoXOZtPS4+yfx9ZwA0rsTQ1BvpBfHCV/iUGfcbjkSrb2/E7MaJeef6P7QHayiVYOzDDk8Nic
1ikaD3kLNV7Tq7lqdiVeRUlm/zpzMW+u2nwknjhElRmtnRn2AnJ1PdpmUC2+0jUSEot2jp3hVF1l
hO2DTylkAkvzNGxuQNnxZeLOhRTgD7jFMGHZTkIs3ExT2eYjolDFLxaJdtMUHdx5PdsWWG1CAJOc
4PP/Osu/oiYXx0ba71PnlSNImEYHV3tzrNA+cTdolAyBYnszuMiJQPoI/mIgIc/g3OoXGQQEO1F5
ODvNFtbpQUD69ae7BLSsU6ds9gpxz17Gm7w3hmYVuvAh5PsSHRqFDxvwo+sd+j2/eMZVIXqIbGEL
9GfQjOFOCd0NpprA5kCGrWJjghbvGbfqCvfmt0GxHbthpMnMEbXkxgV3paDVgM/K+ZOG0GO/K6Ur
Eu0rEYt/XjGGMLdvJ1RhXscKK9CxKFMg0Os7y48Vsi+ts9j9wPapC8NV2t/FaE+zzjXnVg4liHf6
U8eRltPrv6q882fG5R0io5IGf3HsO/9fy5PfXuQ6HWWr7waMbEKK4624sDMSp58m9iqdS1IU2uyn
kooX5q16zt6maqFk3rZRybgD5khUuQwbKmk+DvIuq+nvwwGqzT10MfmD2i6A7W1uku/LwDhGthqB
JTCmfGPKmRTHHU7TuOxG2LFSNOchooPIXKA/MWIAsncfYC2/pwMNgm7mHzugVbMxRUvPIFZ2jR7y
z9IgCRHj12icRV3qPwtQa+nwQM9c2HxRb/xICEYMrq7lSlOoYTWw2hAWU95IJw6XgnLYhwrpcK9A
9ocpZ+p8iEcAwITufoeg+NNCdqLgP5oZcnc4MFTe9ouSTHnrXgDPBaajmYDOlVE4PF8O0w+rDZaa
WbUW/wZy3EDQo6irOakifInzurWmcZGiZ1jqACYs/0cySBp779YhefVjNx6ClkWruAdhWFeY5osV
tzY8AzaaATM2IxTJot5NicZ51mQ4XfVyJgTzoi2lsLKtCyFHVTcELi8zGKO6V0m4hNgse8v+Kcd4
U+0yc+rtLzIzPWuKKcI7d0Bwx4oHYNGIvf7ugdVjCXijE2d6JjgH/9ay2iw84dnJE9HBVrEb2EZC
ySbLJZsQPttgkt7wUcQlN6HAJ1uEsIHHoglh9tpCLxlJdO6GR0lRECydnQbNRmf5e2J5fZaSop0y
T+zsLiRW+Jvxkn6bCN95FSS4/hdhQu9Xc8Qmb+gqdtJ5vV2iPOOTk+caZK4dXqjKBC7nejMUYVmR
ymPFxxiWK1wGuZ3luMLqhyusiD/vsA/z7oSNDMKaODrtgZxI859jW0EmNWA/NcsnZnTPRIS+xR8S
KLdJvrg65mknMDUv5ZY+2Dclrvxj1p1Iy1eHVvBX/nOmHrmzD+e5qNOUaagHM6NiIS53ClPHQ7od
RLNMf1986d7mUcnV1PhN4GDsbJcSsNlgD9pznLH9jP/kqw+POWSdo40rnjzKZZcfjgZcWppxpLTh
ojpwhf8KCw6AX/TmAvZwgPXGdXYDH+1171AatrwU+4WtRriLHWFqQUyosrAo3xmsTAqCUZnNaK4i
BhESCUE8kX7sClejJSVDajHjSTQDlKx5E/MXgCLjTMszGuXqcduwnIy3Ta2ra7DgszBhiVko79yn
i72qcBP8yydDrYlWtd3a+Q1mFpK8tyaqCFf9BPnvb6xHBuBFHzyCO2agygZHA1r2ucHf6EkxBp4k
TqBlF3VVprspCXs6s2BCS/Me0LeEki+Kk3phEnZmuu0+DamRLVYLt7Oc9EMhyXEB89Lsau9agkiq
MvSWHhJjCSEcS4vxMtcrynhoAXwwkfd99xvg5jdc+J/Kmtj0lSmES1pyok0ZOHrOALprkqFkKjOf
7hCZv2OpfujNCtCLEHC+33Ctrp9uyCqg9v0w4XvdNI3Nbw4caRf4XWQHlIEjXwUYcnXrTIBDGOHf
HHFUDEMKZZIpaaPa5HhxGD0FhbITvyiaNdDot6Dm1J0piHYK2x/Az7+SljZxxwACwjinw1JJ88Yl
YDhyZpB4/gCovPs2Rp+wufGyR3Njl9Iu7cYKYds5oChCcJbubZT3DaLNcRRDDZnR03X+TyEML7jg
nNwGdaWbq8b2BjEEKVPROSHe52EmyJN+1xF7WCTvBUdXHHVAghKQuQUH6U1IqDiAIzyZmoPHBugl
cFk6Mm/iSwq3Q++wxDNkay+sSsthDNDyu7N8YdzeEpv4O5tRxbA+LiS7xTDoOZULp3G/1k1FDYm9
Fx1y8rkEwn/sF7Ll4LXf4EAIgE3zzl5QYHAJtaI9QgDx2aVMdvmvqT320Bg2/L5ulBHBk3mKTKi0
Gt+MqPj1mEW11x0poFkqYQm91co9aWWGcWoZDJuTy+HTgGwjK0pG9+ACH6ACsAjmJeacBuIASWlA
6ioUsJdZcNxOu4wluURoDwPxofSQjYGdY6mgH4VU9gJOgRtRSLUzFRkWdlLAJ73/MpIpVi8zDNcR
VwtRK8mYGkP53IxCS8cU1UkVKdjloQspn+SfSPUzieUtAN4yzdnwcu96Q3rHYcw55y8O7pQvo3vz
lrf4pS2xjvHDMvdgUovQwZ1+NQbCMlwzqD8EV/M7JU1PR9lYvYqKe42rosrfzQN61P8DaaR5a4vP
GWkXY1rv0780ZbkbDbsvFWhkmaLPzbLe/chUNOk8qds080DZx4PBBcp2gkIXBD1IM/Jn76EkWlgn
3X5fEzCE1jIhUvxXyhahhEShh4EN5+knTxwWoXi6mJjUKC1GIW+xD7tUrdW2GYrUugkeCN3BarAB
pqKlg0asBfiTa6RXMZhQHKxXHY38WwBC0szi1+TYIMjygseTaFMql+UVS2aKr0mQIhSSZWOyK+L/
/50SRBGhTdW9OaTd9M2Y4w+VB5TcJm7YQUDN7tykbfs5QMDMBJA8XcqsdjT4a0nxG/TJKuNApjNl
56dWlHiDbizbyYdnBMHwQ6vkDy2N63LcXS/1+55yDDQSIEi0bvet50yTRAYo4epArUDgQMscPmNG
bRA7Eoa7HT8X+7HfWFZYXURXFbkzoLESL3aQUrwXs1ni19Qm0yJIXsAnwT6VfAP08jWfvgkI+rAl
R5IbdbnWiPxATABUv1IAtdq7bpNIpky4GKckT1Ji72G1g7+76188BstO9xt9qenmLrmawziqenMg
yqmWtxW4kavRWv2CSSytdT00RuDBD0q/9/eStUI5oll4K3KDP7x6JSZUnO5ZqEgCKZA3jbcX4Opf
7hNj+SlNAl47Ri8zvJYLEGLAqLICwr7qfaSVJdGB2cAJMS2VmRWw5zlCXPh/bazg2rJEbLjfYkjf
MDrpsk1jnGx3CD3uCm/Z/XY2VDunV095Zts91ohKGpeA9RUs2TUdzu4LqwjJihaUXpiibyY8l0Ps
IztqV6/U7JvkrSumVAVMXJEPLgYSXfhBaEOBgiMoulirp4637K8CO34BrQsBgVkAE3jLbYLxFeNz
jgN2rtRj8XkER1vWVwCQokTQ1rFjd9W2i2jY4UMG1HuGafSaxemeYAKRuHXuemIn004pliRr2gyU
v9o5WMJKOTzh35+EBqolDdgAh+bCBnWnU6YoIV3rDF9hKjOdJ8cgzfeW59XY8Af24YD2OtKOyQ6R
mSYF+V0qDrmDEOfIKaTtnnivmh3H/hHlzt4ZcVKLtYVn+1CbDo5B5mgA7HczE4OIkElQZJoLIzag
1+p7orfILrLqAAV7JM2aKoE1FAAfV+ieNgzebm2GvJlfIkvKdT+hLlaLgcMMb6/9A38ZUjXXFzob
7WRZnsXh9HC1qza1U8WnQ+RH8a/1dNgRF3SJRt0cinxqrhE1mURz5Pqjwh2YBjjO8fnZ6WcYBjD1
So/5kk8ikUoNDHFY9Nw/jFNxTInlHHokwL3KEz5sIZTRZ9B0ZdSqQLuADjFf3s8qWJvYKR4V4Nvy
cN48NwiThpWQzZ0PG7AT0A9mKRG32UdYxUcjbnsKAm6HOObcB68zmxp48yY5/6dtHljwUJ21o4K/
yp1EVkgIVonaYjJVnkPHUWnzL7FVHwQ2uP2RMhxfTEt05JQDyUmtqHQzGlP0sRQGVddwQARyHGMA
0IZh6Ft/8Xzy6j9XiOLk2BX/duAxqvLiRshcP9HAt07x0Sd4QJyW79sGH4a4qcAL8FLuH63JN/gp
ZDUL7NjL6RwgPjAjeQTTODwPEyuDFXPNsdSCQFVZcHbIiK+tLXRUTnLVxFqDQ3+DdmU7KigGcshs
YK8U3vU1SQ+W4dCiqYw14cyVnDBWBMZoTdczH8MahqzW4iIAOHw5r6Hyz4+bweeXx9+pTlhMUeTo
JBojhpzB+/+2AnoOLLPxd3soMxK4IPY5VHLkXMDRYcMK/CInrlac0mzk4AI9PmlcXK8IUQgAce57
1jD2PyOrdkRNLz8dYiWfZhOHCo39ReLQ0RoEorN5+m6ih5FrufhJisI61P7pziURdyKnnuB4nc5M
wBHeKR+OcuvEDP2uEPLbxhvdH9nL/jqfvIHOQCchz/KFlIkFg8N/xP8JaVUn+ldz3jkomEsO7OZO
ssFvZewWfR+S1CDJUGil86EfngzXjw5XTUB4m4m9Vp9ZKWoc2TjKd/CU+mfwGPOSR4vVvrYzqRMe
LC16DmH7RP2dOExZbrL0IvJcSgGnlYAIboB0G4gyUHeb5fwRRPoreB50W6huLLydnRdWienqzgH7
cEEGFRzsfOoNvp8Ujs763a2REDikB1IiKzG3HyH2uvhO10LJIDkqBHsb4DmYBpwMQbYe+rftX/A2
5xLDqzZSj+so1/UqGbNAHGXYn7LKtnhNKVToY5x/krzjknJTR8XTxAo86L/b5SFzK2fgetl4/LyB
Hg2dyu+3ppHPWDwTrJboOZqFZanjzbMuoyzxp6B8sM1RX+hkqo6khnHOB2ywv3PL+ZIbKXThfTE+
91jm4R7m13/DyMknuDCz2y/K0rXPb86BFbt1EjNm4Sw97iL2CU8/EBiicSMg6BhQaRLABooFE9WU
2G2eVWRd1NTc9TCruvuF4muovFrytBtsNlGrelpFoFItusZdaUC4Z90qWm673Ja4jBt615o1Kzso
1CyHzhetSgAN0qG0Wv6oFlBTjGlpF1aRJOXeOZLOp8hFV9qYVGEV2bUAvblwV4mR8NQHGlKsppb2
c6/gLjAzT/MZXXw+HqziKXpV8NKW1JiWf6/n5CIGrqvG3P+G4EdKiGISlrEkLtXjZkaGlzqJ9Qz6
R/JQ3Vl7PnNMZc0987jOg0IooAbSI8yjzS3Xb0WD3mZtuQEUOLpp8wdrQ4GzroL93ZDJA5Stn+G3
FO4pStFI68oxzBjOE7WztAreEY4W1bYCN4AHS3utB/8rsSZFZQ+pd+7Jnu45l3NYROO/NOJFm9xg
cCF1lSy0zHluT++UHdTv+VzEWkf/a++iSoNcQKZzh8Xoa5HxXrx2m6x/QOePwNM9p9OQpGV4BadY
Tcue6dey4e73sKuf7nnjR9u2+qtvYeAD6hFTHYIfSGyA8TNFIWZZilfvBS2jwXQcp12aBIt1R5RF
d4mW6/XEWMD2FYRwOsmq/eTWIMDlfdJh/A5UHGgHAnbd3hyFPZFsztNMjQQqGzx+Yc97/HfIfvxz
05vMSBTPadz80PAsSan3w4HoyzUxu0425FH3xa6SLCRdoPMn+xTcquAPMrz7K9s9Frt88XeozVCN
ajM3biHE3ytvW9sT0Svkzg5v7KNMedn+JSadFGct18RkX+1uZCvY1Vq2xdSi6dq+GeONFeNrsRmv
eVM3AcWdI2xPxTvq9VBbbvWYmh9iX3/GoweFzf79EyjJbZR2FjOhoD5/FNwGxc+zM+Zq/SRv7jR+
TQLLU6DOvUTfZUG0brRHKRE1q8oDOoe1xcsjzfeAoc5kggs6kxKFMcn69QrMpnC3U5Wip8Wx9evD
drNBHdIdo2Ag0tuJ1BR8P1MmC8LLS2Fhaoq0gaZ+nAuy9pLJXDHj0f7s+skSq/NlhBAHC3fVcAH6
cGYFee1AnDVIMPzLHIuKUo6E9+VsScRPNUYtw3vqhIayLNVEwKuAQziy2zUucnjChsDx0vsi6xnD
xyC3YFzOzrb9S0Powfs7duARd5/Wa4EfgSsnlV4/fy3yLl2qaTKGzSN3/HymC3N1wFeHZKGVmV6+
Faxj1dOH8VjSQSOJY6cjMG4m5bYh33gBU/YKwFXbLyJ7r9QDD0ciC537veg0PaW0J/InLlKSXNR2
ctKk+tTwAjm/JdivGtfZ4176zboq/PoAQEGURfeF4H1Jb/sedDiYRLvqYXHWS8rQNzBR++BNbQvA
LsOpg71KScNMDrvBjP0eT8izbyFmMdVDqLwNTMuh9cxhazFh9r4eh1G0NYRNy0VA6uZhGFApLNl5
J9J2xyIqgIql7lnBL7+3EWmdWKfmsV9mpEIEUklf1FmNOZILSquvbdw7KkjV7XyRClw6cbauR8Dd
ojX7Q9B3FKnsbsPtW0EaG6Xr3sQ5hzE13fGSiPGS4UMfKNIYdMwUl3EAGMaY/f6M1ty3AFkfqen+
t2DbqG4HByrOOIQaOYDiA1Hzh+4C9BpiHcfFkW6FftowL3s5KNKl+TCdswdofycT3Wf400ifHXFm
gYR46n4V3EI50DKLFfESSvlsOxdrUPklv7l6UfQJdZpjRUnvNygGbxGgCLXhQLb7oucB9IGBe3Rq
t2wK71gDDprH7+KQgcLaLuM3VJRZozef5zgxsVtibs6dTVwzWjrx7cA1uuSFFeczTo3ghZQe5imh
qv/xh/N/Pb066zmEs8xTWZTSSQhaEzzL8DM8wKyrYAe3ZavFCy6FJpcI1TF4DrKE9t6/2oaUHFGS
5dJoNQiR5W+JGzyBn/T8rfP8LRnCiFvc5ClmVsSIkgh6w7WvD/pdj/jDk9BbINeeVy3+Xs6Yuz/O
CJ2MvhFyocGds8Oz01dYf8dffySEpc7xzCDaw9BfZ9JJ2Sji1Z05X3yBsQCxJVmVNu6iXEEQgGWC
3XE5EheaoFQgVo/6ddvvO1E0pt+EwWyFfY43RyU3eYzotowTXFx0EUctanO63QV17YuC3NJiJ1wj
1aTc8+t7FHlepwZITdm441JtrpGTKgItJE9ez4+3TdJTZ5J9I5+CzjqBCbT/AKc4Rq3vidjczHUF
vZbYYyRHbWFhtwqzHX/3mPTUV3I4SIi01VqFwQ6foR2b3HcsbujF2IVoT3rao+RDWeFySXHPdMeU
SZzE2o4+LSl/QKgSuqBtVtoIwP9CLN8RUz4RPavmvnY3OTLW5vNqR0FZBx0CRirkCOd/uhDp96Jk
dCzvsK57cAv0ZPB5fnzEBEzaFvanF3gpVDkXjfP2NC2Fi0t24D1mqpr+4dg3+mtEWmEEzq2yiUGv
4/DA2SuvHsPQAEmltCPG9uBkPP2/sUq6LQwvrpLYrXyu3O8jjVtg0ZjzLtrTqI2x/3EePWodp0My
MZHty316kWXhPwOmXRN5dgEo7O0tTFkTYj0mqVl934qGE2ODxQ0652jxTrAuVAmd999TNT5tgQyq
PXOYWV4qh9rNYJLfRY/KezRFP7ejHFWoQ1thWbeQo1wrlVjXma22Ch7Pqqz+nzsWrLTdpZ4WdE2F
ljQ8LzYRcMc4QCOx4hse1airiIaovNzRPlSPUNCPonoSDkAgVSMFeLPdcsCnA9nflyKZmMtgHCRt
687pu88qrPG8vbtN9kWr3JwwTojbdV0ThXCGcJa7IL5vcBXYP0kZWqbLTnbrqgmiJkI/Md5dwl8J
noctALa9UBufBIbhJb0JTwF5hWlYKuqhM2U7cYQrkN4D/4dxPdSeu+zBpAWITxOJhO2JwPva2i9K
JjtnQiPUdoxhLWxH1hACkGC8cISzdmy1Us0z44EHXHavX259e/Uu17Jwh/8BN8pj86xXY0BaHdDF
pHVjEgyiItC/AortvkIvoCzEsT95VC4zOjBRVutQWtxM4CAT2h3PBpVOhuTQVQ+ox0yPqhl6pex1
NIhF9+PLS9ASExrEJXU64q700PSpxGoynBWWmCJ86dBR82uxCMPbhqNWIu3BfJTE/koqcuCM1k5J
B+Qx1qfbjIYLk75Zyy7k4tEnmVdWo/Rwi8toiEhl0MUt9VM7cgO4gYc2gjmWCGJUZ4jKYGMllD4W
P0dJA3NxROAp+Gt3wlggf4aUZFUC4Hr2keqkwMBG3VRKwYCkaEODNvqpt2mqy6NC+zPXws9WUuX8
PJ/QTAYG5oU12jbJ5n9G4iC2KG9+DrT/yF8jXEPpybQeo6ji5jh9QBjif3ivm+xtfYIOpEK9EniH
vOQkLn+mxaRKrZVQP36575v+AHoYe6Sw+SAESxzLbfL5w8CZrQPGmyfvnJGYrvIbvffQncT/WOuf
KmX8mNqmS+b////CYbXczjarFY1XI04T7VxA804EawTNt+Vdiqsaki5vmIfl4XfYt6UDmAmMz02+
ebXGq/yMsuttuU2NwejjORFWVQ/G7NhiznC0biD2D4xlCana96wNN3g5O5X8SVE2WcBop8w8ytXU
Gcd5yJZWYy/6YXWyDBTbkmO0Vv6zE4URAouJ0cl+u5uK5H9niGsiT+R+taa7nsE2I5nOuHHajqbP
qTAUjStnAyMd36MurD8aQjZZMoPr2F68YrqaNpWOx4ihlrvebQcxZgyVlJC7/pHOwQngYsYbtz+E
kpkMfa5MPRwtMy7LEW89HEmj5ULB+NSrl4oQC/eJ1BnF71OxiE3OAfh6mZds5JJtLztYFrY+aCR9
LmWz4RHIk1Dx4s+VbkE4UlzWJslvTp6CukJC4w0ry1AtXXxU1OC8tDKRnJr3AgREJeNV83ZJrlwk
LRJQDwWCzSgakUfI2BoTIRBylJCxafvgohaUeHM7tgu/Fw5MYrDREi0F8awkmbagYIf/9wTJyMVI
9JgwWE1PpHd3swOrT/fMRqVqb0G1z2Ev1PU0X9NGSCmvcVC++T+lOaqsyhCoAcrjSQIlq3Ngu5fj
pM68EP8ZdenE9CllLWGe7L/S4XBAd96a4ylUOP2SKI03K9z1i0sm7aEazZnuhXZGBTf8DSTSyfsO
3s/QZCNXyC3r5Z0P08ED4CmdHDtRIM2P29NbNfLBfL0/jntyqy9oqHGGpRmvlYh3uzMOVrGzave8
ul6J+8uRG/1FeUhrm9cvaEh12ArjZyv2vOrnxajZO7XOVZNkvah5qxtyb/usF57I/glYABaVLKhX
Po6T2Tk5IFx4q47gKUgy5XG+hrHwSH3CA8Rx1WYMf28WWvtY68XDBCWSgUJqhm0GdCqgPbD8V+nJ
kxA+g7Fc+tXnrjJq2j9BogWDTmWmDOYemWZTn+gVSielZJ8eRicP11JQdOgPJUHAsyBm2tfsHMir
AWO971R5OE+LFSSPKkgq6aL3GO4RAOU+hCNW7rIzxycEUbiJ93OFc/IUBcr/GCHzcCsd2aPANkua
v1zLz+wUVlzy/WWVuC/nvolDo2MkRGoaCXt7wYxQ3WvEoFB09dj8Fmqn/8K0ix5X2uXn/+oxGn4v
DTvYMQplfUg8fmoG82LxuUs3Hq5Mwa6hreBfXwLCNb9vU3t+3vSyJVNAmBh0VruaM2U3pGLa/gnc
7RqeVeTDE/Prn599xDPfj8bpcqERnvEFhs/aU5symWFP3qkqhLht8a4Zp4Zog8w5F+v5YQkmg9Y/
lS++erIfAw8DNOT0jnczO4mEt5pxUFi75Jgpoz3NvpMKRO0S1Mn2H5VPT/qJL8qPvf87E2lni07F
WdmbpQsmWU9ss19z4FwQJwCsfEh+BULsU3G3flKpYC+Mpadu91s+CBVV9Q2dSxjR1KpV9HSmNHzA
y5SYMdeciw1MfDS7c7XieqXXN8xzhfjrZBUwsh6e6FtFA+5B6oJpSFxQzSjBQ2un5Zhn8CldvX44
hU5/0yhPfjkITBz1ECe4rew/r/s1JklORbZF01Ql0M8yfQBdH4E/rkJTgSGXzF67zGbZSvPNASyt
scBvS5SzQ7haa5QGJymET1JVd2+GhMde6SAZosJIirX/aaFQ/7fMLpYcNEkCHWFX1guRYg1mZz9f
UhpozuGiLUi3LTd9drxrb2wzt7lJs+0eojM359rSPQbn5fiKJ/AzqtCX5TFqkrr/aMOSI4Sv5C8V
6obFBpTxjijEuwVUT4kFvJKOG3Tw1rUw3QiMR/b5XyFWyoB7O9vQ/nbDH5gGpsx32u5IQxxVaTJ/
uweK5i3vt+VDZWZhbZgFY0SITGm9qNUZZrSNYgXOY0deEsDDS1IHkaF7t2ad68Ez5WWJ5hgN23p2
1nOF1dKcd5FKnQK5eTWKgbHHwbhk9elh2Aj//G/mR58DpXfbgnHmjuYWX2B17+kiiGT6kqb11OxS
99Hxip/SlSAK2SBTSI3esy5Ud19huy9vQ6tR6LjAPWHWdD7nTQG3WhyTo0lgCMEdxm3iS5Y5LXqy
9vjQFLkSJcFbKLcwxyJeY/TTOJsAROFb28CTu5EAojcbsSFPbWZhFcDmpD8+T8Y6tC34LYkXpxtl
sRHlHOtMmevFi62HUBdJCLgRWr1GZI2andWRuZc9L3gOHIOnSLJbUGAFoMq7PPoJMZyUWtp8CMU2
ZwZxEo8CQ+zZrBSqh2pQtbcq6mPojq1YZVa3UbPS+cdZ8CaveJFYmno5b/lh+IyOLXFUUGU3bpK9
ex3s+dOXtA2O/KviPAscIS49uRxrtGIKRxSd3qJoTZJ2ctInlj167QGod/oAiG5pYn9PaiftZ0os
y3vhrpQa4KnDWbZLzrxnZlfYFVdCRlRoBDF8qhb5jHT8K2tqQbov8CVotGq5YD/pY6WxfURKpLzO
Yao/DKKAPydjI80NB9zTQfS5ESCWIndJbt2sUJtGI2pvRgAa2R7cRJMrrDoadn9et2bKoUXWbErH
HnJPfJRWUoj2Y84KU9Ud8QWgYHjJ7XFoBg91m9rBByq6BLph6Z4SWflZJck1yydGji4VN39SoXbM
hglPs5BGEw5ZStCCAXEwI3rPI7M0h8tYQNz9z7QYpiDUIf+gH2lxFyqzB/eeP5pkKaJiJwva9SKD
VdEkjWhRHRVhxGkf3tvEwISrGcFyVjuyYhHVqy/hT8pJXZRulOFqvF7WQgSQk3UTY/aps2vjJnfK
q6kM8aDbffh8VzlqFB73VTxcf5lqcYKyr0pKo+9dmXeyd8Nfm4ovrw3od2LQfgcB7p6sR2/dSEUb
X1A8GaBEw+f//DIhRVcl8PTwTQiWPzyLspUXZkEZTE8QQPHICoti9YEkJnaQAqAlGkaprz76nPjq
RCLtP1gdxQXhwggt+YbBpTp499uTfw0h6BT2JJKHPHbqa97X+2vSGjXFWtbzdFatlzXRJIVLEB1b
+018EnaUEfA5CkwIQXqD9eCV9ap97NTA9EJ7So12LgrW1oFIwTIWG2OR3Gx4rcSS9s5qaY5Y7ukw
SommpowfT2+Q9RG5z4DgqAHFRvwPDd0K6mTMBwDITLda0HA3z1hzCBH3wLyWYfFOYYMvSDBzR2HW
Wu0WLqeuC21GUt4fJ0Vp4h+F7GRmzGX/hzHxIw8hNLUzl5US2+AngnyP0yeH32bwYfK38QE7OSyU
Jv9L+Bn/E/1UErk+H5oQbXvgeiHSQ2BSOYhHsE00vs7UpQeBAzIfQSuncGp/wXDy9duFMCG+MK2r
a7Ev4uEWl4myBliBSkq3YtCOP85Z3wrz6xfzWSQ2paqQQ4WWsqbHcpzM0T1wXnEl7hOUrun61Cg+
YU/h5RIoPjkrxlPBTHR/pN5AvPstLMgQLwoCL7FaR1vW8XTkGlww3mtLuLvIvuxdKXVJemx5CfPV
1JFaQx0W26g3FWcND68WXcKcw251ZagG4gR9Dful1jqp5JWXwICrNdCkT6E2HcdOnKOrKvNGQHhZ
R/tD551Qk1ILD2jMjaBOqniq1vg+xqj0YC0o8p9UV0VAoNEPu/w0v/qtNcj6+ZVuMjRb1RgDya71
s3wAaxy5OtsXfosybHR08gudLMIevnW1JSGDflaNS8z0ZpFXdyWjGGBrHAYRLrc+pCYapTuLeFcZ
xs22oAtvZ1pMCiW7jItAf+0ZHBcgVwjL7YVUVAPamAZWYyyfSWBb0a7pqXbJ+9aANsPaXDL0mhk6
lFBHWrcYn22a35qkax3R7syVbPDmuIn4twxbhGCd26hyEdVxtZP6UX+1dGeOPija5OI3GhQgE0vN
1MHdxJKyc9JnKl358aDVqd6nC2/5ROP3427K79pioscjk2DUQTEVlomr2osSzSCGMrQ0ajVaZDMx
hreByH/VrratW55apP8+DWBdT1vs6Nl0kYC3lWxXqxK8kH05fvkx/EFmsFhrsDJgs20h+d2J1Shs
6sx4v9wCuBdOyhitezlH/rb7VgeS1Z4lxcw/aDVe+UdjwrpUSSdhObyv5waq2WJyX6bu1D4spoKN
gKkVMSiDXESO8TiXT3lQWXP/4l3lJa1vmy85m4aXAjfbew1engg3MIJiSaBAMOT5jpL0uhLVlx5x
m9RVT1bG+kjBD3h5NoLGYqoe6Byy7nsR2iTdTZlNMr+/so9h5+ME/L4dcANdqTflZLq/gA0LBW5F
dMIA9vpxCM7QdejGSYpPNTtp6UBB3u2KyMjVDiCeCw6GcH1KA7aV2bxnOVQbTR5s/GK/QIAOnIHB
dsTV2YtylLz9K3Ss9Hgzas22CwCbm/dCVoSZ6L3gwcuKq2D9igM2W9Aa0hhTOWHsTUMrc5NaPAE4
M+7vehaq72y897Eybl8bfOcFlq8MH0CHo19Xv1TzExuN6qr5AS+1nG9zXGStqapAEJj9GeOT+KTj
Gx8xRQE/Evge4UcuTs2k6svRNL0ZIC2Cqbi/Hh1YwENp47Gg4ykJ8e6qP5RwfipUMHs5pk1fD2mg
+nw6zN74SxUZC15OOweu1ZQ0sxxY+I8RQBqTrpxPHep/Djc8VXnlKUajRLxvU5hT3cZ0JX72HeL4
rS3zm3GJJTwozD1aJFIPijGGlSvvebufi3o/IEZzNjhZhr5AF8aPl9gZ4Ww8pngtf4W1Fy9nDQbi
15qZfUXiIrp6FJ4XKGlxCo0Ae4FWxDeackuz4A4tJDBl57UUTBuwfLkN/90Cn85ld+8jjVjp0fq3
wko7J+VX1pIq2b6D4EOJiRFhorVtuiTNn2J+Y/xBwHFOOP7ys52KpGd8Mh6hrY5DqUHye5GDcKob
P+zpe1vlfni0Sn1Zi/XQlYNMeWHYdkq6sEHM5drPLe27wRs4Tp453OZl8LyoYpqjyiPhruqxttTt
X4l3/rICRLCQD0Hr0T97p8kveYxd5r1ub+8Snbh0jiOlPpnvmVkYvHFTauAMc5cIhSV/eqU8/Fuw
aoB4vZPz+P67ifNJ2012gFDmF3dtlZGOOIFM5x8Vub8MUxQxwuQF9Xk4Bx1aQvgelhB3XKZ4JifT
8dlTkBQsy3KRidetCUWbxOJqD6s6Ro9EZutNwfW1bzMUN3Lrm6RJ6z/Vy/QCTJxtuThZVm8VscDH
Qq7Zxf7BlkHnKqxUOUiNSGkkPYaKR8erp91cLlJEatydBgjuoZvMVma1hGrT2CKFvx0EPi4tvx2G
UzfiHTmzUUi9P+zIQZCXbtIS5LQQeP3c34nDWUvUznXrZXbLUDeTC3aEEScIqnCUDHbuRMoBh4ZM
qUn0lVsxUER/VXiOu3BkaP7YM3t4z4TfgsPk5Xh4fRpzDcNmJrSkvOgZ1jKoy3WvdB+N2jHmg2eI
INZT3hoXLgdYGliS5RpOFST05cE8pKPy3bwhZeu++jq3iTCZNgxYUrLf5GVnC1sOx4kUDZhm3YSA
lSnNbLtOEqzX1AwilDVE+PSU1LC97s8ecM18yL1YJ7zqJAOFciaE9bFEztlq+OECgRX8OzxO0di3
ZgIXSq5Yl8PWA0XYUEc5DooHw0PdE5eJfjTx4sKfGh6hFM3ZJRCd6M1oyl9ca8ryIDDhNlKqTyqd
1imYZ8/bQ3NlLq189A+xjpnlsHIzFwss/6027ecPGCaQNa5GOBs98GVB5MezapB8L9mOGfiljg+d
9r753L9RVpScZZB+fwemz9ugXwMKsZKgyx917k75PrcLVHKXimg9vNZcM/X1mFV7taB9zUScWu5r
xVE49R06xvLOjjlxSUeK7oJnFA6ogNPCv1ttf0SyG0fApfp7Rg1QKO3AM7Us0V/yVG0sGiCcf20C
CRYnY90erXbFxpLp+HyTQUqdVsr5W9FToLSo/LBcQ3qXU4XgH0+pmPRSu9OLr93BrxLlroc3LV2j
RIXNUG/Mn6z3cTrRsS9wyRf6evyFpqiTbew8OpIC7MrgVgFESf6kKf0fpm2TwA035zk1tqjp3Cgx
QPttlE2QGs0b6PlXuZidJiXNT5AOOD2s0LrEhI1i+nM1dafJvzK7xsyt/2n+H45pQ/C2em71gMUm
/dFWY5nzY3PnXBeND3PdaGVMHIvgqKk6sKrFUS0ZW+OkGkqwkdrgUoBuKpL2luxOXP3GFgWFLC6+
WecmUQ85RByTDCeW00c9ZPYYciTaDg4deuvsCR8HEOetGMRZEhSC8Jh4BPOFCGveKrF62XsKN92h
p4eXiDRHREkvVgdzxMxi7XHKkh1wCH+f/hk+ABARp2EeiqClUBqAJ5phXz5wIM0Bqty5J6z+m7Za
wQlLFevlHhIB1Pu+wpMGi7CH89YHoPRAi0V+dwKgejwQpXkvNGBb7HYjFqrJQhQ7Go3S2pw1HFym
3JGshDxUa+HTchDVSS/lpfAXwqO4LAgHL8tcbI2UZ+I/GO1/lgJH3/rqkRir+lMcJhGv0nFQ76BX
jdvHVyUCMmIhkJhgijgPDa4QT/PbQdj7YisoIlnoiDyeilOAcrLUHDEocsdSN1fg/4WZQApJS2fr
23V1LEYxxf2OWCw4dsRbgmISaM4ggHQo+AzYd9EL30lSja46sXKBKsltYLap0YMFACcCds8DKU1D
BRlCLpNuMOiDx+xU14l2Fd/QoV3BjE/ueTNNJIe6Q5adSqmh9jD1Lk+CkmRURdhV8ls8QFLl9f6T
Ao7SdO1DyqanrfZSdBpTN7RIS81N2aKHcVCHR8uMt2iZX8f/V/WZQhagE67cvs+mifO5/IEqx/tN
PAF/Ph5C+V9fXH7xlksMcskKrZydPUF+hCVSrfztUeorgFieltuhM8GJQaBs3DnnLKHV2xWNm465
cfICcMYI34Uqk42lNXc3jJorxOfnkDkivqhglL8vN5BjmGgWFN9djagQCxUhEaCTyjKvTNGZBGGZ
pSaQ0OjF7Iu///G/AmbDuOcmZN4d7+92ma2P9IvNdNa9BMTC4Qt7EQApQnJlYd5KxcPVFbzMtdJZ
CRU0tIhhtIdMzctsJQOgGx8jqDD8yH6cHrLp3rDeyKh+vucxd6yFa8nhUE83W+veEhuLeSQCIvTY
/EYOYxd5zVgd+oghe/RRCJ09cN1CPpN47s+L4tfoXvW4FfmOmsfjEjjY2HKz7owO/mEbV+Siv1SR
YwPfdUg7125SDH8N5sTSjD9ZQns+Z+20lHAh31KyNPWMusNXBAQ6eRa8pGEdvUgoClk/nCujWdkt
hbnt2xCBIchaJC3TGIm9L3UoAgXZjFdUFvAG2PcSQYrrD18udtgXKYirpmNaM7aPQ2c+euTEZpGz
Rg6AF62BVDVEoU5OgdVdgxjdGBkolT0x3NhHGUDq1i/q8vaktw2Vd8Q5WBWW68lUEogxjp7tD287
KeKGWaTay0YuoKqZOVKqNmv5o66l+OupqIhbsddPa1DOWy9ydE2M4n1yCmZorYl7ZfV3/YspWYhf
UrpjEuv0PKEET2HkrDOFIRn99UOiAOg4P8b3JzaLDGq7P4bZbGFX9OocZK+mRN4nOAnf7/vHsyMZ
kkZj24Glv660m0a6BZw0NUaqYTuBwkNi48oZV5JnTTiYB4kbwonP3mDhAG8jNE0FfmArq6JsUmXg
0DRuPT2iVhz97HbQ5fsmZ2iXvO9b1R8Zhtq1GQQbSWncHsr43YpUELeiwv+TGDgre+EE5zFRS59l
J7FA/YdrwDxpuUtc2eNuSdRRzskzSjafaQYxmy+1D3KLQr9CiPyKeS+6OcsB5dp6tGmdztc4Y7PF
OGE24F6k23w7hMQTfaindqMH0BhBB2P69F3oWFegBUqBCfv5SHUkz1hF/Bfd5n4RJSE8oU+fXVJB
dLGo8QBhHgWD6aQYKMHiuRpfkHsXhO85/z617Varnu4Y8G1CKVGfk3EmwoCTioP0szD63LxTC6fy
O5vhlpfH2F//omhMx4dN4Uw88UuDRja6bU5tLhaCuX4ntdZuem8KQCACjNbYOM6FQepUWk54yn+f
DFK2cSf5+uuXZtOUCLswzAwRSi+AVMy6bskY0ILfUQEhaTK0leCTWCs6fS8NGE4h+p5VkT4iRZQF
iCDEEbFrGhxS8lo+26kg3wet0xa6rCUdSZN30Hk2H4FvfHIA/pJqPLIjb9uVutXmVqZexC10Hxrd
2dEY21HNsf03Ib7FW2WpQrfaTxWWs0py7zir2TMBICw/4nVvt5ViVhel4aucS2bYx8KX9mgLMGTd
u5biv3MdZRIh04ekAEZ9nZa9/U608iaN5hMddSxvMTVNRkBnYE9zG720iGya3cuh7+PZvajPRxck
4TtdxIlRQPZ3ISkvAzkXmSgN3bm4Lb91xCqsngPgTd0ygfIndJZ/QFo6KFViTO0KlzW1THmnij7q
fM9x0K0deZNylQ8COngXJt+2xfZM5Sh6OLzqQxj4HIMFUBwzDCwAyRCxB5u+bD/+JkGb/LMwFwqf
vMqwHV9po0qi4SiPXX+TMQIe1OxfEBgM6IJ/dG89mI59cslyz1g2GvjDaAGbZ1WgAYOSyfRLQ61v
pTNJ7Xyf5yK/Y1O8iYld2ywRBeeViM9gTCwjGnWyWbe5o1i9y+EHNQ8k1FWOqvNJ1E6XcTXn2hqH
ZXa5WLlVqgch3az1LugymYZJTHB8Scb/ovka89npKsDT5OK/qDLA9VAbWyGVnmqPq5xvIc2oi8YP
UaX0cCBnXrSJA9yxuoGVwmtXVGa/pgbZOTytOjgNR9eHfQ3dK/5lP4KHO7OFu2NscyZzhsFr6Nql
Q2uZR6ldckvYTrzyDZ8VxeOvfN2agy3g7y4feY8FYZ+buPg/+lozDlXJAa/M0UHewXLyZSF3k/f8
lZNMAVfUSl6b69O3wAMhRxCDv1AcrqEvHbQiO5JNQygbkN6VJ/5fOBBQs2sudbbaj/Ryo9q2usBe
f7aqx9F/iC/lBfuQl+CjJHq/o4Us355g+z76MoZAkIZvwW6OhuN/jwG/FEgbHvWaHVaAhzTEqN9b
+JRPONDG8/4qHhrbiIBBFBHgR+lS9IV/YLVe24njokh2wHtGvDtASLA7RSTsXZmGHnmeu7AwTyZi
R7I1nVki/dMwKIyKE3UZrNuJmfDx8RjXuzQMfG3RgL0Hb2dUK1AYMaLdoyOzQeytJndwOsYcX6aW
Hd49psti6lhPElL+0/fbK7Q1fe7qAj/6IzJafHUucmcdMg8N5yKJ/84ufItOhjTpPDUvfonewgdF
e7oMpnDD1pSZJxywPxbXJ03J4lJFZaUTZQPGwYPMB0tXH9kMHieZK7u/tzpVwTOZ7a5C8hGmBwMf
knZblTu1CVKF5scSIUNVuGQNorTG/xnJJtaP306A/9NtVJjYK4V7Z15QEwmdwderAVj0qU7sOedw
hVVt53DQvPp3bfQy6GvW3ITSz8+ej1tO1XiXn+kLmesvTlTAR1j7EN2mNGJHbqfGlevQ64pPkIBF
hkKVZeWVVxHb2ZDZGCsGL2pib1R8By3eUNqRCljdYL7l8PDPU9B5q1PBE0Q0pUKsUIDQ0eOcuD/h
wnCfsrd2aNf5cYkNlVYYU5kSlOZxHm7a+z8A6Lig8P39vcPe6X6bS0Nsjtnxgby/pzxKdW7ZmcZn
tokFqW1RTARVCoRjNXbC7CW34bye6dXfG39y2lCH/Xd6V1vRf7Ie0x2Wm8/uyaO1t8imDahjJ1oo
QgcBUA8hW8374Uaj3HPWk1JAT6J0RMlUXt7uaEWb/N6ExgirvKNgYtP1VbQH6RUCjPH/D82aLEMM
j2mNuHLI0Xn/KbZmfJPnizOAIlc3sl4IsxU0ukp2AqT8pO1oIM1cxd4jZ35tPWkauhr6XFkyMImA
QyEKp/O3g+5Xvk9qT9a//+kkpC3FePPQXLPeYgaVJj7q0XrMgI9TCJNyCh/1I/lm6hHJHKuj7h8p
LjaaAlpYvJvYk32+BPcHaCSVgLBQbb2JkCiyZKwqLi8LY9YuyPhJuXDFk/g/LEzuTL7SaQrkSSKd
LnfvyXmbABTWQzKQsF2LMKhr+yQTtSzHe/Bf12VWG1hmqDui5pB2TcLPpTLJ7ystWRPGtdoyUnwi
O3Bjb2qqCrSi2FAUWDtCD2Mw9DtNsyBqjQvhwSKC3w4IaxQMQBzoYAx9V4LmPAnwfAog8wFTAqBR
uNp58RgAzNOynimMeaCjfqHNpnnxvNjIyCKQx9pKkHpBcq6EAD6uY7eNT8JbcxmJyOIo9lNIA77V
xOWie/+9aTWZl2RUxWLPa9F9CtheNZ4Tt7Wro0JpkDMSezeTameQ2zOob+3rUR5LBlF7idH0yz7D
wpdFeM9aAUchtYdUHdsjgae8Es2F6P2QRTsqYGHXPiGvkXHWuhFhtDp8LVybsWoFg3j8+tC2AFGE
hsY5TCDpyC+176yZ88Q+rr9gmi4lA1TVi0JlihiSRKZQw4/zwc1lDblGAvkUQEkos1NYny5ExE4O
weFjv0w0UM2RDw7EOl7z6pnCN0GqInO6UofFai7ZO2To66zFRMTsutHfp6+gOnh1p+0bstLykpso
73rwaxLUXh97ewcso7ZkmedZTHuRjQMDEVEoTYC4FoNaG1tK0qanqseljV1fjjs79QlQrqUVz/w/
RY7fhcgdBU1XR9AkAu9dHsXKgwIPcQbyd7u1ajYwJtpriwZKUVC57Gw0BRYMwAhEMAqJsxsZcRLI
WSoOtzYpyatPEWvOhqPADIOS907r0he+eM/L9APomHqNArwVNsA4wqs/2Dbou7oC22PpuH/2EbnV
eufZPwsnkD5kk87I5PHZlt3jhSqhsRRprErKoZiQXg97Rxlh2PZyyuioyFDyOyue/N2A/BW4DDUk
bVSd3b1AKPRygZ5+KgkR2cHgDAuEp1Jzql9+kRXShsRxdu3CIF57r6ky1+QbmHZ909iNRICwtl6Q
9j7v8mDu0t4dN9fRDaBZRynOzDNYUAPkZR5DHf42CGnUTd97QZmkGsCQ57MK98D1sQYbGniSHOOW
D07JCVZtlx1L6b+/OBNd0Lul5ociVFR2JJFP+NtlpevdRBZ3+spNX5WeCknenubNysdfy87elVLB
tcDcc6yOerqdepudxCwXwevL0uTisko+W0VIOITvPeGwAuM7VS5QdMzgcV9ploWSFAjXX1J2Y5aH
qWXLTzz8BoQbE8pjJXIYBxLpwIIrsA9DH7Y+MNtVASHmtqX4bixVed6Pok5FsvdyG42ST12vH+Pd
OPUwaTcHdUYY2qlVod44IiPpHn+5waBPIOM5KTxN94ag2VyVSGaCWHe/mCmaNPIJHOnSIzOYdvhT
+pyoj8xwnhY7jG3PGzmb7Mg6BC5u/6kKPWbDhBoMpWX2hju1V7FsW33oOnF2vdVv9sZ+YKgRMlx6
W8QBWGHNm9qWetTHhGsuEvRKBCE1poMHJAYoUaW74OKOQV+3m6FUcLGyxZp0m1+H6MCZQkGd0qRc
aFV90fofIQFqnNEmhkmZy9+h44GTLW2SBFMCx8WZcucYQHcGHft0Vbu8TakK4UUZtHrh4ENfuR6o
JgwR5B6hdiPqwhyLElJ8wP0OcRQhkq+xXBZS4GVuKmsSg55Dl09fqNCrXJwWGl7pTbMuHY0mff0z
3Kas3ikTzDvjk4VRPQ/L4HIl28w1pfCOFDq7FDUhSYCp9MJt/yvWzayzvCLIOh788S6aFimYjo9B
y+tCawiEeMIlmBAA1bcwK32WpAz8gmQqx6bX5U001FkOooCk5fc3dwR7DgDVmYfRwWd+HHNxKsmQ
eG/GbKCPB5hpI/2Mtso9+QqchT5WTx3zD25Od8WMPH7aE8jWvpvc2F3EMW719xhbjXEFoSbj1bVp
nHtX1ZEvshxzZYdyB7Hl+QUPtHk5eN+aJHtPhllDbJP3NyADQKE3IpNY0paGTx79yFP/CYQyxk/V
qLoI9Ecbx5IorMyzV98RoNdNGpMtKEdSvocBb1AuU7co8x0re9nOwegpHF0eCGtc42B4UpEpoVEw
jUWsXjJiQqT2/Rt9Vi+PpfjuVoQWT6pwnQluyHEGWToTCQj/NE3GR7O/9q/2Hif5yPbiyXkSWhK6
20ETVMN0VOD2XcoexRCycw6MiKKn4yrsPXKSc3kwxCmaya6eDKepfWHrBsiwIDgXZM15IzI8PWSf
q1fXfdrWfomkL9ZD1xea2JXCeSZVwWImcLiOxB52t+5ZpegYcyghyxJLOCIWCpFBtKD7rzaAyIL8
quwEujOGDI3DbKYvCucxwGCH+1kQu8XSMPBMWx/sZFHhHo6MuWGKSHAiMOHIgMfMJ2qZfIsTfP95
89PGhJuIQsJ5cQg25078+j8b9O7O5H21Q/fsfX7th6SR3ER7se2qyBOxMX1MKsInPHwuVnZLtdbV
HBPqqaV45Ic8ONEI1gCV7lINNY2yVJKNCYWJKiCLcRrS4pmrDAFjMi4ZlckKSvUHexXZzlN45aKj
QTlr3AcjYQKnCfGX8/iPwtPa+ot5+llE93FRD5bWts1q9gjHppCYQQJ9U5MWPoUD0y2iMlJcFMED
awZN6KHsVseM63RfaMDGWzIzcjp06H/mwbhpfV6cZicbMni0ZlmpDexOLECGyWxJdxU4pG4kMo8W
jINZcn/NQr8uIASYUh9hlJySCur8TkJEE9ouxqId5GKnDmmQe6Whgns35t9h2tjPmQLXe4ecW8+9
VAiXaXAloQ0rdZgOvjFQ9r9i/wPyK/wurIUGetvoJrIFRGSi9Kb/VAHvQA7pniC5B5wGseCyN+z6
3q0f60f/5LVJid6sBMTFSUjFln13pnf/fxVo24hTfMYB5bn+dyMhJvaD8pyNa2E6/AR2W2Wx9IxJ
kzPP5afxIrfWtB/7jpSSNAGgrVjPLymqknFZCXfawclRfwUsBDu6mba++vBlywW55Y/YIw+KDyhn
nDYbR9/lV1m0oua8xo1caK+jMVJae6CYAMK9SnESRyc7VVhV06KUZPb58B4YMWGq/74P4jeJhduU
0H7LklOC4LJyGKC6mHmS+4cQLgYt37SMCGRL5LsjLGtJG3vrtHlh7SHwe/bueKDTsdEXx134vvoF
l5+n2KMhuSFI1aHdxMmfqI8xn9Ib8nslI5NPkiI2ZsLa9v58YqBu8YmWw5avk+R1ptWcnV1x4QQo
hT9l2wXUIPTmF8HZNOyAfxR+iF0CE64BC4XPqZXM3iNts+JQhiG8I377cUbAYWZtcBQaMqYIiuhx
phEtiN+NV8tPCD0kjSrcKPSCDbnB+Yd0qVbpHA+zK3IsJfFUwBsZ7kjedU9tKD55hEGzO/erdIAf
motFp1kCq5ImHRfqTOpF3711XOOs/ko/pzH+Hqhd8KYAPRSH054udwCOd/nFx9h8hf6AhJowZbu0
vL+IOFoC3co8nAbZ2Er1g8xVgmXRtMDEh9goZQ8qftt6M1KXnj8zqtuAW88+fsHkA8UDrlNLXSzw
V5R/cUA/0Su31phw5C9cHxFBVvek94bUlcGvtr/7Ja/0USd2gmbhRbo7p4rAoY/nIaf2/jLG67e/
XfLxROa70jIneh7r8tzirwY/RTjlHfcMT5H8PNMjeCa14uZCHtgYQhzMjffZu50Bf7RbVKpHPeX9
w6TdAwcer0sT4B7xSvGjkveBRXH8gQtT9OSemmYO4koOckpTB/MPyOe63OgM3Sa+1+BEllhtVCzb
2gJOKzTSc0yb/k5dafFmMWW/MvPWWLa+Uu8QsHtB4VUzzQDAt4fzZewgfFoFE4BXLopbOnXRm0RA
+U2wp64QJIYIjtLH1TXs8oTE8oE+4xSsMkqGYHljixk0akPkUTLsb4zOmgSTljMbTQVIkJpxqiDk
KqoN4LLIQsqemi5AzEn6EoERuCIbaM//UWkVyfAd+CdIIA7Ba9rtjfXFbdMhvHlSdU6Zn8wB9YqS
CbgI+NjnDhGYwqxrvey+ec1aKttp5RFTD326Qokv4aIhdGKKoBRzkJbFrXhbsWl2FE49+usoAfbI
kL3CJ6Cld/3qTQI0QJHm8zFp5nVYM/gmNZdjrgVvQpnL6EtKI/y2X6czTXPXnuwLKZZ7xHb44KxT
Uaw2BsG18XOfR0Bqjk3jVSMeOVT5osRcbvfrgbDJ1It3OWdtC8ZkEBAnkpefh9SibXfe6gGmJXqJ
mWj0tEHwISyZnktCsovscOI3lVcZ4+7Y4FkzcKUXQTWWIZhuRnSNFVq1jO36qYo3VVb1p76fZApa
jeoGVba/iHnqwZKuRkKXSt+BJ2flSVZaP4JMtmQ7lJiBmvDKDsOkcQLQO0DVqinFY+Fr4TIH3xbn
P8Vwz5b1j17pwGP1kXdZtjz+N304mfv8W+7PAlavcj2FvZREd2evgjvYzYJjsokff6uHizLhm4RQ
zaTtrdUp3I+9nYjcPNOctfhzRzY3/Twk/5jbd0zucxVncQ13q9r5mResGdqr40ZDM3OReS3v8eNz
e931lDCVhkMk2NwIYyvR16iMDlY5FNNsb8C3WE3t9kuVUyqG3rqIei5CO2kBYmUbEybK4dAl1yhM
pXrFy6iqtne+XjwxC4ObM3bmtqvFjN8cN/dvLMLjZwTSI7It6XnnvnsZRapW/wJA2Z2BZ91Lb+FX
EWwFfYZNQ6DV8aQQqoEJ+AkDN5r9Is0N5r0Fn/ErkGXpz2NFcN0QBKiCWq4MuSR/GDwMUR1xiaxu
mFAUXFFoSqlYG31x/b6dKlPNNQr6rHfxaqJDEsGWjnx4TNZMeZCEXaz4Dr13bt+pmemNgeG3E1oj
ZiKkrLBWs2VFLizCgbIU2jazPZofMUFCeG6vTvYT7Qoksc5+BuxQesLYjbwLl3/ndVkPuuJmW2vH
Z0ZarzbjXi+0Oak6S3AM+GmjgoHif8LH7ySL0LQLh+6X1k0GGLB8d6Vk2hOZ+WelPadHlD2/gxt5
Cn3blu0cv5OakMZj1cMEM6lSTbhh+soPRK63oBdzFlcQMqs0bne0NQADPk48s7vI2r4wRd9eVzSW
1nhNlUr+n3wL4rb2qcEyW2GqvWFUhOpL+ybciuGmLKIvRkGwLG3nFjg8Nzd0bZy5y9lhxWfzjj06
ILICuPa+F7JfrY4v2w6ah68qOTpMPP66c276J+Uc0WBEgVfArBJpcwTy/xN7rJ6KGu8Oc9W3Ss+5
d4Czs+QkX7INeYGBJUDMjIDMmeBPkVV10yFoFZx6tr1kNJlWzQKCcF9yJk7rr9KbXoelVAUFLREW
vEVJN0KVstH8UXeJPp24em0jR446gp+TlVtaB/26Swkg3eXH90ttiHxu4rfdnBHY+MaafDkv/jXv
yXFMf5/fA8IJJflxEOoCuRnKvCvqpod1WOa+12hXyeQcyJ7yMnMaKhTdbqaj6Q836pdArevQUzTB
R7ybrBg3UMYSzTZ6oaRYxWCn5LtZias+tAftLbPnsmlggE+xB2/MuyoHW8HFN49L+4jd2rfgB2EN
DQCWsExVZnTGd0EVB0pTy95KHxaJ/YZhFAiMluQ/RH7yK+3I92LXADjJ045MOpqPHC5wu78Mt1UR
gQbG2Zd5rIVl/iC1iKG3yKZVkaCZJG4FdRk/Czt7pmgKn2OZQ5+7hIY7xYmkp+qM1sZQD4fYr2tI
XoWVR3rjwV2aGIx1zRfo+OnptLAMxmicsibMTwj7g9XUFFAVW81thjJ53d0dvm2RQEja2kMyouTB
hVUxH1dvFI3cbrUqrz6GacXFZ4Gn5xQXUU9FjWP7ff8IDw5NFwaW9jEi3dwk5LFHw6XUnTG27MEg
Y+DdhyZJt0GaLrgCyLO/M7z/8wb3vuBQGAj3D7aOjAIgcq3jFBnXcMEKVDdYkY9N7gmCeRUFPnPz
0AwxL2xImGaZqbTYm+1xULJ/JisE8FG2y/RwKvBRa8VzX/qwopvYX3IIsNlpEeBTNRNO+RcmWgCH
Wc5wG+hoaAnnBcsKK01+kQEkl6LTrHiwM3PEt8tJA45U4at1C0OcYESIMN2mLSimWmdRO62JHN9S
OAtsRm8mu41uTKjFzTOPM073BVMiIbB1ipyKf6x7g+bLbCoaQmxqYJjpLRJcfmpBcpIVQAwQNyUh
ONABfoFeJ6ZDRj0t0qXIqMU8rPSjcuHmi1QbbRbmB3qHRpXJJXNUrOsyT6+WxL5EgsyQNFAjy/Ht
BVtrl9I4KLmVjjhftNuO+e3AprC/hIrVTAmC22I5vAVS0CYVmMXSMikeO7wBJ5N08NHTYmmQRy0G
JLJ69LXwXujlapRh0zdiOfEx7QQkqvedgAZVb1sRlE849Q9OHIVyqlbXgYBAdExhG4F9ORAkoIMs
sSMqhb6WClvfMSr3BdqpPcrfS9Z7emGywLCkXBH4e8dMnyf+sX5XSpecr2iRnl5ZKLWx2yvSpPpy
AFOTbExV0fZlW2eCIkpq3ckRiZUXbBVUPw7+9gQNpRzi2ROCPTTwPhExqAms56xnBMl4a/rATt0d
r2H8cUUxE4XDiz6PzEOyRO/KBB81lrcAW0MUfphg+EHrJUkrZgAW9z1+yddl9oFcv/LEnG3Yt7Ll
hl2jiWqEy2oO0K2C9i6AzbNP/kaeF9lbRg/Qq0XKVLAehMn/9x3t/jSUI1iT30NB0/1QQoeYjIkK
Xgy1JJeNuRJ8wQTONXJVfqehxSTILvbMM0hMswT3G05qRJ9rPJvY2QpK2DiQKV/ACztcMyN5+WYp
DeuT9GO9OOEaSLoEqt39jh+XovhK2UdUvUIVlP6FVTMCPiugctqfg8F8wVQcpoR2lFuekt19dHMy
PzpU9rvN9+C6mhGUs5+yHwtm/NPYuIBWZwsJRyCV6eBgzr0KH48wFOSmsepQYcW00mC5uNM37HHu
l968Cpl7MCywqZataaWpaXKsWdz0wc5xa2P7/pWimhYorNJxdVUPDij0LfvxKOI753mvrhEGCE2B
FhB07GtAmq5ETuQ481mz87rO/OI5USlwzREf91PKYdjdB/YK+RjdYCQt0+hJaa/IncV+tII0Q3K8
ZMWxw62fWIukJjfjCR4A+8qbFKd4We+X6W6R1nBKhpTwztTgnphb2ff2zjqN3/r76+297QeFKatv
x4dH95N/9AEBZBspEH8AfE0lkSTpj5MQ+HvufYkyFye4ZRqizCHXZOdCgbkf2QikdX3Wnsewvjbx
ZRyH48grBDRxY7OIi30r9dKC2YrJUEoLXo7FHQsW4HBKD2AN/gQgSkQE5BBNiqBCr+UZGoHvNwjN
3rHqph09+uxX9PAnAv5gfledccrJACvbiDHui56jfh2g4iGB4h0T1CFJ44pwEUZf6HMZ+AugBOvk
lSIbvA6aoUT4Ojg/PwNKzlxynIbSA7vUv92/UM+etO+IOq5BqUpFTcXO7NakQcfU/ULthoyheR84
f6TOqbQQz9xowoqPA1k6dWPVPUFO0bKaGI9+7/QAR/sujJ4eBPM0im0korpUwdQqmw0m4ySn65Dc
xa934Sb/kbmN0Rjk1Uztk7FfHPIw9rT5UD7O24cS+BZoFdkv/s2fJS2Sb8/vcfs9p7QYPzYiktkT
WSICIDHsZLO0GYtWh3yVvZULUydcHvi+SgJkH7WoN8WeCmIruiDzWkMuSVyopYM4KTUeYq+mDxuX
De3+JKwvyVfCxMKyruxiO/JM+r6PXNEyW52sH9SS5fegAKGC+zRWb8BkWWi7H+oC5/X4WQwurwAI
NmdWbPg8yJYqJPLukrzzbpuGp8DDtKxh6+hd9iqfEH1gNIaqFuHqVWHuM+IjkFR5Xqv9pUde8d8Z
yajWy3/EeSmBPv/wOKhE2pQOnr5gtZRISpgh/GhC8U91WZOZgUsRjbm85uJDtRuzop8qeliHAxLS
PWiTk8iQngV+z8NOzuKq8KGsjt/kCi3gaoFvRpK5XXjw38Af/qPqJ+cTbd+//k/LWd2abbVYTrbf
jK4prEVEtX9W4OhOenWpaSGBnQ8JKWU/DZEraipjiYj6/pBGUH0JxgjEm8cSNaV7PY5EczTG1/Eq
2CAri+YVktDZu7FMAO2Q1BNclfyEJk8+VJAqv1z23gO7lPh26N99usJvai+I8tG4WktIMAXKIYFF
JPrM8jNljmtucWvZube33lcmw/msvhI9h01KPjjfPQDiHPQ7QuWseqlUlLCxgeVWqkvkO4Tdu8r1
zgU/14EDMszFtv2LwRn3kAqqmHdNho13TZpJAbNVz8Kmugut6xMLUCHNggWJE902U0ZXxqKKlLEW
OPfzxpWAjH843I2aqJ+LMst2DV5Hi/TEvrtawkqeo7QK8EoSAYzfm8NcmKHZsNRWkXF5lU8GnMts
W4fXxbackZx5VQbacV9P03i7DDVTGxpqchMbFiT2jjXTxxOWnNzlUCoMH9KJLP3Cg8H5So9GuuUX
v2IN+qt7zqMIj1BlWuKkP4yv9sWLcbmPY/VEM75Z8a7tcafPeFMAxU8l6Kymni5J3tlJ3GIAffwD
4Gl/FS0Ymboi1mmj/gkaQ9lucVBnl8q5vPw8UjqoAbCWB52ObIlmu8lsobYe6Ts1IP/jttPNEsIs
Fsd1FgNw8vCWQdq/VYB9t6TnksOIUGgOUz3ElEEWRgsZTV+aAO25l1hbbR5U0ipdNljhfRcPXYhe
znkyQgRh7Uq5V7UQ34CDQsNdJm6q7qvprpxnH3suiQJhDep4/IFw9vqkntIfqiJInh199ddBHa32
5JxZ1RJTcsQN5oY7CqsP/XpMstId6XZoYS/k5wopmxigWFaHCfUP0oWi8nAEF7zBs+gVYTZ/A7pg
XKVsY+VWSVfAjCgjztttx8GwkQw48yGP2DBrkj6iChq6dqSlmXAMEFjVKbrByPap22lne9oUfNzX
LO90NPfrQLUGKwucNDH9JbKhIqEggBusUk6i8nqEX9LCmnavj1OBrximcDmcUeVtU9oTaFeBfYzi
tFxZZEahCXBk7lN/VkuHHfmYJW+HOCDADcHZo6+9FBBH4UYdPJ2kNvrDcpa1ZqeAyNjBYBjvqDnh
o7a0sQC7L3FtkhC4SLWLPrZng3rsNpAdN21gMaDCYDGU0wmvJTZRJU1cqBHUh0xF1pctC8fvgWaF
fXYig7DMCExIW+NXEdz7ITGfhC7yijVtKcW9NjMlKwS8b4wNMJn8clbg1zCzDRBRh5v+0Uua61Kq
7FkstZ0UNYIHasCp6Rlqaf+VmYqaBx+vukmJ7j2S1bZEaeLlQXbHZOY+JEzeXybBFikA+cpdInpw
5irSMZfEl6BrgtCQtF7MeesOa1WS7oFPbAz58d2kXZSOsIBRg/rw5SlOA0KUIfyrDaLLgJc75+BQ
13mGSO0xDFynZ7++dQsh5Q19Weg12NTJtdmWzmJuXTsgb8WpNCU3JUD/i3TQgAoAw7jX7+EMYTqr
O6OZB6QODIj0+Ac9s9ym0v+VCGIumiTlJBbkZj+elqSGb6g1GBsG43+xcFLZYPNEVivDhWRLT6OB
NfNhCGydzGc8NPKw8u3L7T/P4L2uunmRZs8cZIMep7VM0kaUyMQmWiPKdvVBEaqU1yL7d2M2CWjo
BSY6COIv+zW4FGGZaOj6Dj4496BR1Af7VyUCoMhq6vfdMT5m8PIGny49ufzHBaCClLk5Fa/o85ls
D+y5mZI15TIGJhLk0SkntW5+pt8F8z/7smvVCmMnVgwL3tz8opt+9FaZGlfYmHYHXgOsAa/1UjMb
f7kR2S33IU6GjrueNov5c4oHnh8p8CZgrQQln8qTUbdIgDVg9iCAAIy3z7NGpTnCxCIDmtTVhbzi
XUlMvsavkaarvoNIJ8zdN/BcRDYsQg3RwFo6ePv4rklWqw+IM9JaDahLvnS8mhYdQLNnWoKvQlsA
O1HxmDNezmOO19WKefLjCrvzGL4RzC7DuJ48SM+eh5Dls8kNhyrTFIZs7+Ea2cE/uNFDCFfufj4B
sPbUR/hRaa0oWpk1P4Uf1BnAtYN4D9dSlpkNp0p3AuIBpA+fnh310xUaLXRuTkf9GmT1Gfo1+g7Q
gPxytNsnsF/4rx//ZQ3dEeGxyZRP3HLFStIfeot6q97Tm/ZShA3ZCrSlKtYFm0r0oeHBiObCNtTr
C7oCJmVo2v7972m4An3YTKCK5N4EfDnwvpXTcHo3ty6gtCzMI98pCVrC1gQ/dkfKDS4mBkOROwbU
WdPbLPv9iVha9IF6AMEgrKrCVOi9wvQRg/DfQ28nJ/+j6uWAQREby/n4OV+IufhcqyfivSlQN5AT
qCODCTd4UWQDxhniibruGtlNcBz7qvQJrXi2jtuPq7iiZn9ORLJYcQ/guEBtnmh1uyr+jIP0/Y8X
gboBZqsrjArsbBGxzjc2QRJTivSYyyuqnv35q+vcFb0dXR3ZxxtkgVRgzEBSDnicF2NnWd+F3Q4J
M9IHKHi2o31QVlM9pkIvWzA4IC/iTWJBRkw8JV9rjormUHaJs2GF08I3+1Lnh44xdh1qfV8FRX+J
zPmhYMYpXNl6EOJqZLdUX7lTl9IcZi3l0bc7YNz/lrnjFUNjpfw14j6Fe5lrN0VB67rhQBgDq/qJ
+/Uv/EJ6h60iLxKztyQT793Yqft0cHQEgLgnuPP+PnNGjsA/kcku0CfqNi3xH9tptO/kw9nfTN8J
88rIkOVbsksF1DXSQFqiSZ2LHktMvaQflalKEViDNM2QbTKzA6bBmKLkNTJDmv77Ciee0ZgiIyt3
yWg5WzcFYxwL2W8n4GueiXFOP9FJTazaNS2DlMmpZpp5cO20vDv0tlKx+uX35Prql9jMMVVLAcxO
ZHQ9c9l1rKGJTenb3GXNsLn/4wNAPYM7AsObHEqNH+mGbRFfqJ2ay4TSVnkRNkW/FalwGqa+nq8n
rL1QWwzzK4BhvmaLiVUGVyDCbgbV8a4WimN4slf47rF5swFxxtczxvOGAhV3beVEUJkswv/GV1UM
R5eMI5+mnq466wbvD+Lg1RMpL5wWeU5dsB+oyx4e5RWnjFqM+Ed3P/ZP6sBg2tr7dU4UV7Q2QvPk
jiOX3mUoLQuiVWDjQvxxhWVRbJk/LkWuanB6KxAVFDdf1ZPTV9EyURocZ0RVQmJkMVLrdTrukZLl
ImgV9NBFFoYE1CpiVPA/r6a4toFpb3pzW9oI3XZJ57dLddO7AQ7Vxnc3zWYUGfJezjQpCcBQ+I2C
sMnI5s/FjOIJbRqSF0ouDg6LOSwJnq8e1IVVAuP3EzNXPevAy1VkOQC+8gJUcXbmccYQdJX5ncLX
SJT0XSQ0wBLT5p34rVEh2767lwTx476s7lb63+bn0aUJ/N9YXTlUZy8FR03m31HWGrombuk9+Kf7
o/1bLNJxixsSuYBaLn7+lQAifXh5jPwoVBGaqTF99wlxHJyZYsco4UxfY4FfQqrT2yzNHaqofGVS
J0aq0XzWzj0B/gQCssKwIqpmLj92+iZk+e46vr05M5ZSna7mz9kDClkRIfO2XE3keSTUg59Cz6Jn
y9jJNOALdoUFI7jvGmu6Z56EcIQhV+wbcAl+0Mc6KVZvSenqojjm+r4Tdv5pYv6sDI50ZxZeqc/5
HJwaWVDQcVJwOF8acA/PP47R8XGgNtIIw8oahd+aPgMgO4HvdMz6N8PJ7kukK8rm3KrOmds1pG6f
3zOTRlmlFZvASeIbPolQHe9G5upnLqx3uGryZyZHuY7aocslbaOjvX/YN/nd6SPON2mOG1nKMOla
lQpulV5m/ZW6dBu3cAOxx7ZHl97vL5dJApZzaj/vAg7p2msjAOKuthzyvTj5nFkBotr3nyUw47WC
Q7CXRwUHJNPltcJGs2VPOOmBtmzKYUUPMMlTC1oJF9l4LlVZpvxH1VFt4pl8U75pu4B/ZJz5v1e0
rT4TcEzdGZrFEK5Egw3J0POoUWDgcMLnsp4xHJU0So/hy7/seWdwYSnVpwNmJaeVZu0f+W9INXSx
HmkVNx3/cZwr1hnZjsqn9c2xqpZE/VhpHzYuYmMvqAMTGxrcVt5Y6URItUfXg/g6i/43yh/c9iXg
V3IK6VFT5t+atOiR3g5mZfR9BLer5aHji5vgKjIbSj2rv2GypfgLWWTMEvB8hREsrYfBbYB5DVad
vsmbes37QSj6Arfv7eppI7ycKeN/r6Ep0ukrXdc/5JAw8TFsDDv3octungtJ3T32UNDpPJEmcn3N
BMFqPxzfTezoF3fs2eV0V4r3srgjt1Dwrobmjl1895JG39oGZBVOn+F8r5Rte0Xjy5iGqp6B7uzZ
4r++AHbdkkcdQoO3uddGMLUDxad4+oNxnsKc6wBsqdlmIA2LMyGq5gYXigTz8MnrUd6nPF964Stc
S06rBHG0aXN4vu0AIJ8lQgfpBVm0NVOTxxss9Xa4SpIJxR/xEJQhuNiK77BaYRJMgmwlk2RQ7YHE
M3ir563hzo2dfJlyFcFiHuEDOHK0XYPqgb/w6x28OzDZFeY+aa5ZCcWhq10ZVpUA+LpRiDbHD3Jo
x1VBP8NJ68//YgN3PDXkb7h8dNbtbBgu5Fh2OMqTS+gM+HibE68vo4T/ihihwaJb1KQKX9BtfpcB
hwzON02nnMmo6zwj5S2UmHOHXO8v8NA3vTpexxj0xSVvmwZQr0oUGIMHVOBGYWzdFea/1EnnT3y7
S3fOpybkzEGVgwBub5C/qPPbqO8Fx5T3cRTJUKQDz2Fcy9+n43yTnmPPlQdgvjO5MdRXme+8zKTH
XJktXTq2tkAETxtZv7CZDb67hMkvoj4d2qZijHA2PNMx6m/WsJgCXvkSk3peXT3mgXylOzNCOpKO
weE3Wy0Elzc9shQLP9Ng+3lK4LjweCttOsqg+V+zGWm4NCA8OSsLhRKqPgK31e83m3Qcns7TW9kN
4f+UxMZ9GBhpGd8JhaJqKWU59UaRl76FCDoJz4KA2wAkSfDz/J+j4dHzBeqGGxYyaYBBvonGikUB
yFxWYtub6ZdIDnQeniyhXwBBu7obOJyO6Gi4QGi8Gm8TZ+3FKNglahdUfc9CumSYhG+cdNlstnBv
j5/ZQrmgguerzi9gFokW/bnyJsnuAich40fPMMXrV9TtJ8ReMmTjTfkVK5dhDNIASTKp+43qz/ig
YMwhNRPNznfY7MekMP3iKkHn9VOz0irVXEYU9ubln03QGvdIt7bbFcAAPgvt9AzHUZeVf1mUabB0
JJDvhEyc+1roBu7NIaNlnLZ0jtqh6VaIiuprN4+b7DlybJCqdf+xAf6l54dEOfQlSeD40kBpkDyU
lOfi8lweT5vDP+bXbyh6YejewvTuvsPt5CD72mjtKt9YXbDd3FYA0F80hRTyrF/7bUKL+ghC9Bz3
PakAsW6ztirnakDBd1SgW/UCSSbsPOQeeXmvRT4Mh0VTWQZIRGDuzZkam7cVp7iUwvoI/jc+9hBl
tZD0gYgYFXICA/LGnigpF3ZrVB0pHaXLjmm1UGFpnMf72hV3NjeYwK/9hLzsTg1ZWkjekno4aItD
NmNjKGhs/NFhQPQxYICjBSHv4l83TWtPZZP6SzbTcCAAVOcqCEmPFXVUYQ+AUQ19hDMYGe38Mllu
V7hRy6Y/GphOtgzTVrklrchxWcVmd7tO+by8pxfylExSr+i88rLsiE/eq/Xg4e5+YFwfNWVwFbtE
0Lqza7vmL9yf6zuEE76ri6m8ejs+NfNI1Y2BuZfUp7GzR3XaARAiR6rSEWpdWiWz3Nxglu1rVTo2
rodrCW1H2Qz0gffd+EcMUgkmklIAM3N6tg6jR7vbxWEb8b9gBW0y8GQs40DOTVTqhdijrxHiaiss
vk0hWBYZxRaAN7Qmmw03eMUY0clP2WqmBWwS7W3CLaNW27r5WEgWrHbCfcq+R7wbgjT36j5+F7Jk
BVhmU45UjN3+oQXytUWyISnoU3iyghk2gL5EILE0tuh9cLAtq6/TXxU0V3xNv4wylJlONiJ6euUO
ZzYBlrgypbdj2LuqKHAwU/x4p6aO8Duu2yYyJVEgeTaxv2Yv2pn0BzVVu2QL3zBpMspzvrFMSx8w
Sy/mW+CuElccu4581OqRPCmtJi86eb+hmUa3amYtWgLdxWjTBpYG/6xqByG+0EfCDXOFR3YU8sGR
J7shtYPuOgXizblkUCikTFggD4+fnAM2uwroKCV60mi2tKK3T2Ie/y9Tf6a1crsC0yZQt/7nfCs0
08RuYPK3Ge3+cByp1M5m2FJoOX1q+CGUCFBOmmZX5YM1TFVb7Fad97LAfGCURtRwKKxOWF5+fAXc
FH+Rv9duonMM6W9JIrzlIeowZNU7r20fvWNB/+rBE+gWs+lN1R3KVwo7h0jkDvtZnjDgbyl5ROqp
/qyryhKsZ3O2N+APhy+WeTjP5ibMzvMoKUMTv2dtoqdFymgyv9zKAsCyn0qhDKMKkHEcyO7362gH
0LB7n12ePGPY0/oLGixsyjnWDvaqhSZvOHrlap9wrSVyCQLA6NYJn9vpxXO5bniOSnYJUZfLe/8P
M/717qk/os1DpLmpaoOo9LE8uKYW7aE5rjotnZ0RYoPJoFAnOrEF0HDJqSwHXkgI6uGm1TLeDe7M
rwzPzneECcURhpavrgyNqI5KBbTnyJbmVbleUBi4Bg0AkQy/PADbM3CKZ04mH74YVgSvGujeGjve
Db4zI5KLmjJY3GLzUYUfW1Z9Wm56LWTXoVhmd9tIwrW71qoiJ/K8v1XYmS7TBnJjPx2du8HowTwr
2q+xs9fzmn9F2XhuhXSaKIRiH5vO+zNSs7yRXkU08/732/d0+pZIRmXalC3K9usD6AxwgPDQchLJ
8auMplJlUf/y47Ve4TlsbijIvRiEUQzbT4ACqH11i5Rm9OdXD4tnTLtmKMzWehgQivnHNbUTrRKR
5OO8/BoDhWFkaKGGHPFm7oy8XhWBWMLEDymPhSi23zngkdejjMykYbnWNCKpMXQTxvSvU1grLhWm
vh7udxdWS6YboA+GN5HyoGUr4xTQAVb/fsQXzPHpOCl/l3jOgEAcMaurdqeH0SxaqKv24kNxb8RV
SCpDOM4t+PCdjopb7GchIMfpr2Vp6b0P1d6bqGMEX0jS1JGhEPUDKnvrgr7R1X7OYkztPP3dO2vz
kEM38V/BIAyMIYRcw8ez/c9TveqkZn1mMuJPsx73HyYqaqWC4V5PEQo7DpfH+euzXQotPXRVRg/R
HSJ6tAUNxk3W6YhEqTxmNf0nYipyvlvfQnLrrBss0ufZDvdxzsUJP5hGp/T+Fv+asXBhs0fZg9uQ
03Xs3kJCTovhqWhsk+xfThH2oFJjQpOHF7ctgcBFw9ExmQDaW6DHeJL408/+GeeB5fcHpmlTm7mV
Hr1NZeFg2g4nAMFoMv9fOBerG/ct2uXjvg7tLIxIQN2LDRA9hnT8c2u4HBy9M95qYnTAj1Z8k4H3
hDdxsHUYvZ3eW0F723RYV9exG0++Gfkp6FbCJjwSp8mCwguxYn5ikNIG9l75pW+Syl2lWwOs3Cis
2D6f+bQy+U02oX1Et4s85hQTH3P6Gc2aopkFkF+6EiTzViPaAuGSIxlphJ0rFC0aNtf5x5f37OKK
9ulYgr8SyoxyJFUvqA8QH+7JMdSEqrdGF2FWWIdATY7edoZxLbE0gOyunI+WLjI+gUJDgnr2BgFv
IM+EXcVixcyOQIywQiIPer7DOFynmisDzujFOBpDaDv82pl1mBeVzLzYj3ERHIiBEFhm118FAhU6
LV/jMAPCCt8HXWP84VmdVDnPAyiTDtHOeAW8S08HFExMq3Nal18f4oEioImoX+/6hiIksBj9LaY9
U4hiRT833FqKiFFFdxuZ+AejjFERuZcMP4FqRRRans4K8EdETlvdlR0Uj3ZoX+cvqBNFnELiKzq+
ACUSz/usugeYuak1+Fv0GFiqBPFBIot53xosQ74rAa+7WJZRq5Jhky8Y1kT9y7i0qoAGTjuOoZvX
usIF0KXo6+q5mLHI2iiJiwPmF+unmMu0XGJ5om0EkUmgqEBHWaSa/qSm2xeqimtjvRLjy4HVdA26
00AIqYJazoCNafc8RhjLQ4YvD4HWFgRQ4bst0HPki21cHWnCl9v7NwjN/XUIZdS34abNECjduVnE
Lt5xqRV9T0ElHyzkQLNNG8Obj/WGkg6ssrUQUZCC3hzSB1wIfIM9PW03qI5zUbsm45X/0oJ/AL6N
6rk8rqwLtuFye0KRrecVkgy99tWBu5+Hw/qj2YQP7zabStpsqlzD08OMUAaKoRa40U3JAkM2Yls/
aam9IUXAZMx+CI7Gv/vYC8C8m4uCZTF8KUt9QpPr3FVeSvnpItuyXLz8S6peOXOQ9p7bcQ107ISM
20GM1DmMsi6P7MN2Qcly8BcswgrkSRr7UiMiFuB4aNF06cuZIgVXEitA2r2azrU90ggynxqNvmzT
76/ra6dYolnxWYib+2YyaUGdsaF4pKCvajKwTJY+2joH8ka34FmUzHbwu9Cx7ICedEX/MhKS6DzL
HgH7tVhKSu7n5GHRlxUpgxzapmZog6xziXCY7xeXgPOC+KU8qc1sQXOGpr8joX9dHBffC2rbg0yT
CTvHj53qxPQKfPZojQnImFjVdby/RzqEQ79Mop5R+l7qnzjyWO403LkEPF+g+9Oxw5IoIiFc84E5
eh6dTN0KKUD8lbapmJooVR9zUYwlHOS9fVR5J+CTVdwoof575Xu7UJG0PvsMrOtMFH2FNFkEl/UG
KVbBFCpMW8UdNVu+zVxKmkiGv1RWJ4MabZd59LR9TFOMdu8NFHpAv3O6oVC5jrUassOEJFu27Di/
svxbR+mqpdI82dM0dSZNm0bbjeLryqdXQrGmU3A0Qia9UcGRo3+TOif+bpElAJGwNnoi1Q5IQvni
MX4T7M6YlCV407vZulrfZpgcNqhTIssEz1vpdo0kB4Is1FhmyLAL3jNei/qnFjEUyoUAQlHhLE3I
UKH4ceXPi6XoOT2uVccSE10K+N3swJg/lc+ZGYqoHIXiur2fdoeU67JWn9f97NcRyjs90V7N8hq0
Ox8f5Rf36cQ5tsXelpNGs/HDldwBfqx8ILYSMuxSrdMW+pDTPDfW1qiBYBPzhjCTeiNfZOYm6TdE
prVBudUUQW4qrbpCIi0b51qfa18TWlc/qkUTz3wj+KaFtTIkq6cEwIEgXuwF93YC4MovGP+XrEiP
8evbxZV+MdjMhngEFO051mES/QfFh41f4/vnNHIiECLuJrNh7BJxsToXqAjgpBmk3mvFuP2dkaza
bEHnh6oAaFJnjjHu3exn6CbKoCbvOKo2AfyY7Nf3+r0JdzlJM630s2GWLfsUGR+oYvVfDRCJ3a3L
g2nB6Q/bzo9pUYILE3t7LqIbGmNFM1R9rbVs4MzNnfekyXkgrw8cz7rwKEUbdJ52WBjQooOUFtTu
L1S71MAmn9S0VBmkaMw+2KoeAc8r9Y2FxCBfk7/BHsynCS5rL4tcvJg+6yK0s1YC6P9gO06oHuxX
iIgTTgVhmO44qumoRs6O4NX0SULEXHqWz5avnY4UnkZfyS54DmDc/AWTtLEG37x1LUFcF72VuS+d
I3yChnN9UsBB7SvAsfTiknHpmIhNOeyDkQRlOPG9lvGVgaeKEmKjqTC5MPFQxX+0dW/dUfrEl+NH
QZVr6LJaSWiNdgLhAfKC7HFeHfMZgbkhKXapESWHeeNrRIQd0M0RqkvPrrGmozHFTnj+FjoQ+xmY
jf40EOBG1wVfoLxOPuVGz1abBsnLCmmeS5NAbffjxKQ0B3YXMb9JMFWlcMBhvP5leFDxxuhOryXh
lMR6Ks/W3P7w5saPv+iH1wARRbX8+aP5+tLGaBvcM4JEbwNG6wU2aozbKLW2hslvb8GTEjuy2EdT
yv3QtbPo73/hh++TKmsO7M4oO1eEytsc6sDQAgPUkjMiES8nfCdFXJh6LieBELoori164aLFmJLo
c3U+XD600iwZ74IxxVLPcALV14aftzJwOz/UMrFY9R5l/1XFIGG/HUhNrUo0uwCmwfFD+7RiA3fi
gSxtJeJR8fy+vLztYk4jCorhbUlaONlVv02dwrdoKA8UTMQl1q6b48gRST/KxeGOAP2gJpdIUpjt
T/efG2qbbz0iOuhCxS1tM1dcmK0xGC07gQQ3ckpjvBcSavx6LQKdGs1ot5PsOsluDtk1m2vqaz3S
slA7AWB8w5sEcgc+zNbkm7OXbMDeCGLh8Aj8ilvBErGsw1mpVyayqzAMlQ8pgAgALgKWly5yFTI3
YqfGHcsX6k4XNC9f/8dFOruZkbFaSh+7VRCqs99NufEsl9jsC5VWX7q8bnNVLtcnhcrerv6hiNK/
dhY5izWQEdqpo/mZ3Laly8vht7qbwMUbVyfw9/qW8su9rN8Ie/OC/Ga2qJWM92iZsxzRkZ/8lQDB
wkNHMgKj9beGlCOoH9fYh1ODyoHbXLw6qnnp0ixzjfqB1zRYMHUsr2bZj76f9GPeofhTgAwAW6WW
KbXxFsRrj34TGxD9Djh0htTITm1zhkAxh8kgKwAFGYE6WvwokAjhhDInwrSFr9q3/DwgLh4C5nzR
/wB1xow/j8c85rlamjCUrB6I0ki2VET/c+AnAXdUOKz9aiaox/u5zFcPbkS2NxGFb0zYeC7TR9gv
BHPJWHqw/PapC/mUAyBKYgHGgmwN0wJ5HQirXNwX6siLJWShETFG5r8q1fECTeKefiqIg9evqQhc
9mGIG7O9qelNeNyXxXrKSboOeskCSFasMNT0EnnMGvKfUZEH/fBpH8P6XtXLSA2sSO1+4TRYv6+v
2qfaJCDPu7rrrnrezuTw8EaFQMiYA42uS9rMJskD/VXw8KR3sBOIPG4CcdzHnptPO/FKWaODBnkT
eIQY6h26ivQte99VHeY2bnsQGFv+/WIalLXObyKccTW+s0IH+iKErRAhzYc85JSnnFW8soKvzFGP
SXkgxZmiUBeCphz72IUMSQcYkOmjbZ8iFrhN4dpv5y+a3vcqdFZVUS9Mpjs/wJLbTyL7Wtciq/8e
4Atf+dEt2fGap36V7Q0OpavZXxD9fMG/hZ3dU4j7IrkDjmHI2lpzqxMYVp2inVqLEnmBIHrVp/xW
OjPuCpPzyMUQgG2JkrWfzylvyMCuG5uln3lXl3MTFEPmIjdyG4E7zqTWWPOaggcJr7TFW4nU6ToZ
Ijtu0S17GcLP3fO06AXgMzDyS0Q6LBOWgZlZrcpOpCUieeW/7SHKQcSZcbtFRlORW75L5g/igLT3
mpuxhd9KZjXMqFrKuY5Y4YifUxtVnzoUPPUwSrl+z9Jh845IZyzbbgXC3mbdRN7WZdpypL2Tlaef
IuL2RaAVNYc7E079rrOEfn9r4+9hVXFbR5e3dSV7G0K8pxvC80i5Qd4XroYAfZ5yLSN01JuskyDg
Wdx/A27ktrt4lirvEILCtbY9IFORJyAjKEY4o32FZFvIdKQakpjt9KzYbw2/khCK/gLwqOLvUZHV
LZncTLMaj4sw9ImY1SWkY/prldTfIFR6rz3Fl2GVr62ns5BZCWjcDsnOmOGwXMSEqnQmJLp4c8W9
tFwhefjQgJOgRLEC2OMbXf9nQ3PC+AXP6YWlNu4rX390aE4OV/byJaEP9wo8U+EhUcs4PmynvO/0
Jri8CIiESd+R2Jca3bUI2ok42X0L2YUTfNosSoJmHcqY/EDpIHC1LYnCp0Wm88ZKWnmKrEiyg1S2
5+SXcWUpJY/HYAQ2XBCm60emmnxm/rC+AoVV5pYumsS13IyCpNQWKGYkNBQ85PvpXJLp0rBYj9qw
mlmSpWZ2S7DTpJHvmC0q77uZIz1JVXXfEF2A65WU0j/oY3TGoR1yQ9e1yAFD+kiaa8iJr2l5XHml
L9uvivgO3jXtrPjE6IrzlXZN4CQlX2Tbp5UFLbHtHAt3YqAl1/KQ2NiQ5uscFqJyFYHcSq54m9eB
Ge8g0pzb2dNp6yzbAkunpf6Gwot3UhyWUfXfs7xSWB3/ESB3t+/DRy+v0wEi7KTHhxVoNwUQ7X87
Ft+aOCcLLWXp6XmO701uItQ+shQ1KAhQslOxg/pB7AdUA4viHkTEumLcwNmX2bXCRrvyS/NthIQT
CRHeKIHBukHiRLsZ8T1spxlykTU8ff3qEu/qV8E5AEpFnLxvFFJy9575FG7hbGMjWWXPOdfuZKGG
8Y2HdscQKeC1plQxS/YqikIEVfBGZfAn6KgIQlmogHpPHclqx4May6Vydkq6Sczocn6SSuYtRsxA
ZUrDyH+Bh/qyMZayLNvwLdyd4SpuH1X4W20zZFj+p3GamL8pNfKzm05XucMg0KJYXsT99yn/UmYv
qvDVysDwRZlTJONsoCaR52JS98qEgfUC7xKprqdSGXcYwL1BaWRzf/d6atImq74LKpsslaZJT+71
a7XgDFAIm5zpKHatdI25nMbYaHJGsyRe5szknIHqofofomik8xVtgKG9aJOoxkBtTWwOeky8citX
7GlKmOEZWTiIvuicmGpSrbDLQnWWPhQk/4NAC7mWDjLAd3d7mrquciGDflG1qNyWSd95aZVLjVvb
oH4w0rgyesUD6/huSUGNqETPUARDv0AyqQKsUl4WjTfLUxSHdaeR9OrYtMXkVQwUokgOZXKdKZ5V
qxh8iRMIdq1L1cD+zK5SLIL6K4AUb10tvOPO1eBk1ZO9dmEV6b4UUpS6lf0ERpPZtOrRaYR/m0m2
Cr6WUTPIr/WH7DqdRYGdGdYlZcDQDi+GOzoKsEPvXrX53dmAHflDN70Hci0TXH9fOEcNP2OxH6pV
wqvviMI8KG15gfQ8fRJWDS9ulIlNLZFxmFqYCoNM5PVVKTuUBEYfuMXkvjoynkW9Q8vL2w/B9s8c
x6Bc2hYIvBOGoaSU9ivAwlWOfZ0t3dPEzUtsoy4tXUKADOmMVHJisUH+zBy4KOhNiuOcP5KkHZ03
lnR+1fRyMYiJJLgvh7lT2rnF2fOT1BkshPiqPfCRte+nraFdrs0mEp5K8MGsBhqXbjyFeHEGuxo2
IHMG4+g2aPHPuKUlBKcQm9rI0cL8QtK43EO9gSTBj3veOODPvowNjmfry6EkHtjfpX9LjFCBM0mX
PYjYsWBv621qYT8tDGCDz5cYgmOA2dBX4jnXw53E15G6nfTVikub9B45hHkANjeitKAPgwbs7zJa
KAraqI/LULM9pdgF2rL15kJ+XXJOcWwOmrzEB1j9+lYMA8thgLGCPLjQR1bIZp/bJT3x7IJjOlY1
KSNCmqvmgBhX7dPsfiYVgOSt7UZcF7capMHBPoQSoOWR2rRkIYjay4DyYaBYeITp3KR8dBQ41roD
2XPkjr6FHbO1Du4gsWlqib2ThRSTg+hHvr4P8G4KtlAeIqFDGpbajGwEQe7aFbMOe4/mtpzBiK/5
cPhPQkt/zuG74wydZmCchVcTzUQx0O1pgv5WN+9OB395UTl9rs5yKVokdv4w2zLyKvbEuW0CLQg4
mhuBCdujPEeh8Vcvkb/Y6l/+KVkRStOA9XNuyi/MaanQgLX7CXQUoWKqIaPA6zg9GnznKtuAoYU9
vzP/+lIbb5TIR5O8P2oG0jQYl6o4eRtSQOx91ruonTvMubHyMb9/m/MmosgDeIsDarPF08SHUha+
mXX2S8DXThpbyaEz0hXLZmsfmxuQRH40YVRxiMk6e/OczycpUtdB62b6CFBmjGUfCWlUweDKID7l
JXNWEOj17XXUpMj2081PtZhsr+dIwOeM1bJHB71NTIZRHI+3hfKt7GIZ9DqmVCQwGMpuXUrzXabF
RbnQ0ELyF6rpsT4RXBzJA1ry0W2v9u3iflrAxj+yfn5g2a9qpKkcG390htK9CLLkDPMXop37xmZ0
dA6tPRr8B0bSNNt3GyjfbBJualOlR9d63808wBZ6NBpHC73kahaWy5hwr6ITc/+Uhm9JnQ0AXurx
m1+uDsBTzdiq0XIG5X8rRLlUjtEPrOKnmxgQl5r6qeXPSiUa/EtC0l20UhaeKYkXvNzBlauFoxCJ
CznyOM1t3eFSB20qe9t3aFrWPDjzl25RqcIj3wl8oi6mVXHM9tzMf0AUnldQ492i40n22tr66ZGJ
D16dS2Y9UMApXh47aVXKfUUjrrhJ0icMR99VHyEMIqTG2cpseyH3cxeGsuhdVHEMAiIHr6C7+fid
bH5Mp+oFnE1UkG4Uf+POjEFHGBVfQzSDIQ1EZ/BymZsMld9etW+zFbqLLCTTpL2zq4evu2LXgi+u
qqcCLVkvcCq6dqnrQ6BMB17ndNR6puH9fhL2tLRX7fuUXi0EvLJzR2VUtteTKCe9gyg11CBmcJl0
x+axZD/HYgDXew2WzwIyKR4zHtrr3GhisrUhcr6Z0syebHY2ywCUmABR0GJjEIR6QEih0icKvgh9
FNsLX5e3JA8LN4aV7eKn0H7fEPV9nDlawQ1XV9UtZCProWKq9CPgNenIHcLYLbL9cill/oU3g03c
bFw9+WuVanlUOjqAoBlYTm3mCbk1Qlmi8WvGdFrWlFjKSJWOL8YtdJHFbfvlHyYr5hCyDwIuIW/E
eP8XKqkgyJ3Ae+zrRvymXgJ87tipzhyDwA90PvJRN0LN9hf4YbQRYad1hHoduTN2xzBSPQVRqv1A
vsQbvSotfpyN6SxIM48QXB/fTKcPq5xrZzueZ/79++DI1i0rFSBh70Wb0ysVPVmjy8ORi4T8K4b4
PXiU18Ah8vX7Xl/ARJ5cFXumIgTXezutF7uFJ7Cp5kF71tN5/yR9kOlcivEr59T2McB5l4aEqanZ
aFy7b8QoShCgnvDHZZk+ab5awzlmCV4Eer+yKdvxwZmdTA5GdK2swQjsJ8dLpbn2PhtK8HUepwJt
1Ddpar3wdbDE7ojb5Ti7vEsWfrban6VotKaBtiM3HRJSLQMZ609Fg08ixnHPJZkHqOGkDjvudi+Z
XM0Y4uyIvATvg5cDcdvH6HwyZYg9FXLe983VqpI2gmJGcX51iaGtcZCilW7XOYW1Rr6Du1r8ERYq
CETtgq3LwXj3E0vSOkEhzAvP6mBKG6UIjkk8q8elktuPU1EkNmp/s61e7fVwCb5NUrMZNkq2cxBS
3aaQGP0u7VDRACGXE5qR7+HFi+pNunXjncSga1GTVpYDD6rce8TGcCJWzH1MgQzzdUPlOgENOrEP
e0hH1obYVDAJZ5PPaWt9tvUg43IoM7IcyGVYwt6L5sTG83Q5VRdhPR6PESptfQiuARcvvpECFaR7
/8XTOXB2EKOSUJEQcuepjAXrzbqhruTngyk5s6D9kn4qp9CEr0xAMRh9i6tzah2Gq53A1XCrxSWS
aYJvP3q0CIZyP6YXj1Yc4/yU1oLX6dIAjFYZD/eEt56sJrVFbN1ruRe7kc72DnqSBFnbQQKznrhq
fwzTw48/axRsnTzwaIWEcDovhVZbLLJtJNldNXCravh06vCx8cNRE5EvYGL5Es4Y/jpHxs7K+ymh
XKqEbiX0njzG7Cs8heDWAQRQAPzTXkLQtyVV8GmJ+tbr9PYXoGxBEWzscS2FCBhFJydRdrwiAbje
+jB4j3CFe0cpk6PQPZhx3N95MfEnQSbEX/uamPvbuwb1uvtNuYkSbv8dOUbJBq3Hux20Cgfn1EP0
/+pLGOKB5gE2FvLXRw3p9ZNWO7y5422NH18lJNemNw48SK2E1tJIopsEVB/0KMJJeaqv4Z05S6fH
gKD7Ig98jptftiG7DXlARe4oI3jSWTSnBBzGAIcYoj52HjW/lI80uCEpWQhIiYZYTKS1LoOD3BpY
hFMYvIZ/SQiCjeUXDdZ43YXaI+hifr42qxz0jzhetK0cwvEOlPiyd9tNd+kSEV3dGeDLpu7E8+Gp
sQsG03n7MHQO5QTcQlvjr/bbBzv7nXYXJnyIuy2GEMCfQ8w0FQH3AbJqjwYwQZhW9FemPOIOFOvr
8tW10uwf5As8YUG/A+vt/6b+2jd3KCZq//L9e/XSz+Ur5x3/V4pzTv73i4lBCEBGo7+gGpU7XPGn
QZ82shoIcjx8SWSVoQXJIdWKZOH+8sgCsho1Qe1Xo7f+nDQb1Y4BmaaS+391EGe8i8yTpact6nmu
3USSajxJ1aGuRGXigzv/y7kKEM0YEYAYLfslIAviWnTN84vg0OF9OD7P72Xw/OJFExVjgHkB9iFB
77fO60irNxy7+cPYywuGyxHBbF3okVP1iPiRt1io93FCIFH5YLGSOSVMMts6JSu35R3N/JihvaSL
0OYYuFFj1k0Bzi/UFLGcXgMWIMcqh0MQYTNsKygpA14yBpOtsrgiqavV+7HXVVkN9pU1Zo9ckV6G
1dtoB+z6HlwLsubbhGVwQGVWXQfOtAKrl1lCnV78h+AhVZ+Ksc4p691u81rvs2spbkKctEXRRrmJ
dUPWvwosg7YTY7rPXWDlB0EeQ66noWbA+0XErNeExHqJzRtHY3HsFnErKgFxk8Ziud8GeKn3viHp
XFXB/5Pzvh2CUCUS593GOFvKgr2oJl0orCmMy2TkJB25nqqWH/eT1T/Oro1r9ZRylc/3Cei4nszh
/2MzSOEKQCshk0sbbfiBZ0Yat3Aj9MqGl1nBkZyp4V2vgWSpAI4iJlyy7FNKeomr7lBT9JHZ2F75
EwoIQUoDkbskmoeEGLHLkgj6icHGg84CIsM0AuuySDkAtxJ69IZObCbjv7M+3mvd2kg0Pf2Zv20Z
PVuqLnu/Q47WNMUknpRsvesH31lrx0Lf0td7lgRlOEpo+Zmup/RGfFeW523agjX/foDfF15Ka9TY
h8AKUkY5+XEXkEMaArV2spRrzoIjYR4i3kyrMzzMuOFdDEeaC+QMS7NmA2nd4xyv89MwKUq/IsGf
rCU5xSEF3e0ZoqhYjz+1HiYcX0OeOPzPDygB6VsCw9ggUN7jNvRdPnW+myzTGTKKPWnJMWJeq8Ew
/hTnNWcK51bnVrk+HD8Vgbi8GzpfqoW4DkKiGhbozMzIDtdwFcyeqfhreEKqdmZHgnSIP1ujNWoe
NkK3gUV96IzQXpmvAF+paX4Z+EZaAYwxTRzK+/HoCQTQ35+hwm0uiGJQjH/vDuLHAg6ZbB2fg/7B
kCsKlEu1HGVqLRsTl+SlKsyeKRsUj6V1yP0cEoyO5QdSz3ar7iPh07I+x3xXvA9FVBk2kt13puK0
Y7UT+JXHgxAxLqc/atAHKpGW6Nf+RrpsXs4cYUKkYh5QXVSxeiRUXpygdUbhphXLB69pCc08R6Qf
8GR3sQibJo//deSfl2GlorEjHgv863xh2tYVWESe89HIFCcWPMDqQ5+s/yhqcxyCKYwnJvdPLAlS
Beh93wjrKw7EZiXwSjq5BmNs2UJQdJ4H6QuShMSTgvO36wKpXLGVPQTnsSbK3tcxpk2DdiOSCbUI
ZW1oO2jr6OoOFcXPIePd6VGHvgwe1We6UDG13CUydMRmGUUO+XPq9FojckKpT5TKL3qoq8B65Vnp
vG8I19YokLOxobR9a4a85FGItTtZFo1PkgriVPXaVdB78tYCvHjRNrdIFmuGPh6tyHzW+a6WhRgH
xz3GEsy4wWLGssFESZ14G2vyxJvrDcfh0bCai6OQ459FoVHd3fKDxFFlnxbH/PI5mVA8rcCB/99I
0/l2pdWrXpnKfImzMcKD/yJF6XNS5i1H8THAPLkMBA4zbQgjCyvzBFKJOYFtAVS1LjQJvhhdKO/j
Pp525tT/7ym7bKtuyempYZ10hjdTLRsHe3+2jfiOwu8DW5850GtDLKBYJOZCnS/5TqmWHqW1/f7L
htX884jq+IM0hgat+hKCYssQLoQwK+7cuONPrgTNDf9SEWnjep786ts2OTdpV3P5pDh2qcWoZc6N
eItmvoPfcizA7pnkMLM3sAz9KlC8YHmjjRM2Xz9tOTj6IYN6j0GnHXjdQDw8gAMA1f2aDfIGPCKI
il/MB1nSWP03ACJYL0APVunrW3bzUuN6B6ilWZTmyBPz3PDq/ZXQEGb0GIQ9sNcnJSmxKJ99hfhl
/IzkrMw6Ter4VeBIb5hoI0ymTTw2rid/vCXM3n1ekWdfEle0dBIyY0UL6UG8cfS32EndCbCmP9k3
QxB7DFsEicJ47aTpmvvt9bU940Vfl6F7Fe35CxavYEN8bmljaLJshR2X1MrBfuPFt9TO9f5ptCz5
+/G8O1A4jQb9DuFyPALmPikSSG/j1gxM3VoLnkQ6n2+sbj50AqtsYRgdWVILF+m/yqjf/BsSDxCg
kKYe+ekUheMO9eE3tWf9LyuiM3960hS6BPJT6qtvG8QUA9YYx5ET+gDZ9Dg89yQzahax1z9pJ8s5
ef74VY97ndGNvlqmOX8Mz/tYNMx0urU8Ryg76xVXsVej4ag/OjG9v07fi9f5VsVPXvde33rneUBU
WOV1pML40FVerk81lgFkAKOSa4c6Muz+LKSjvhsXBAIlG8Csy43y5y5T3RVjB5onbaZaQXcz1CpE
DGgazoygVrOLoX+mJvTjz1/Y+7CGlqae45+eQ/49MDISlOZfozTmOInYYwoSw7I+pIVi46Xn52FR
5c68RyGEHC2Osg7mULl9Ip6RMICuaCEs0HNIT+Q035vv9334IiCHSnqKsX0FfzgY6Sf6fFoWTq2Y
4v5dnAbavshFwQtg8N1JgNwAyPH50zZG7c5+GP9Q0b2RVaXFBh7Jh3gF4SvLr5EhSdaBaX5f/Nrd
MinrDGLCqNXRAOR5kZ+OWO5+qyyqe+9Bp5RXGMTGd7JcI8ZtKtyY4GY6kE0DEd7i1QJPLAss3TR6
04sP+AtpTFqwCjrdohpZfzXV+faXd1EhMSN1V5/OvMF8ye83rUFfR7ESFD+KT8AUbxuCpw0PlsZt
2+hKh7f/20zEcokSIgbMpc7eAc3k+DAE4S7k1d67WsqdabmyTwelitYPDTwdusZBCZrmYR+GM1Se
2cJVHwGeSZ0dTSp+Si8K+uwEyhiUxA+61sdvde+8nGZNit6PsAJJR/H11khv/24bivUH2vYwulIF
v3zNNB0Iq9k37fn2qqMKAOFvhHZpHfOM53JcSE5jDI4t2lC4vX9IMWIaP23IVPextKvtuE8qK0h9
yh076UW1sl6mO/+/nFpQ0Sb2UYq29Vt0IiWg/lXDUWTC3ZfDWev4TbRFeVLp2KcO+Tp76AgbDfbj
yubjlzeBmYIbxhBgNk7pas1iEFq/iOmAsHO1ymyF2oeL1ta0vX4VUuuhPQhC0is4nDBzoTj0zV+i
Z4OUW2HRmXhz26MdksLptOYtUolMVYrGH5vCitTKzCnsgtjbXBGbTNOsTnb4YuJbUFD0XkCHCCpC
4jm7MN7VrqWGMXHN9DSQFokYuMF+8OAvy30DjCar+IAD6PCOxGSi33FW3nsle9qqG/vajOu3MMBP
nU+/2XGH1pgF3tCY5jg4cA4ehnC6PlV4Iql7CMzc1mmMGv3IwV0luKV2Y7N4CVKMHQ8rgUjxctFI
JfiLcV22wkYla9tKRLNGU3UeDR1VMMlO8MlqrqzeFiuGTmX24WtsLjvBcRPTpBUNAEh4P1l/YRfS
XeoBtHLpYme7mo7UxeUVuvWN2EIzrXztbloKmJXzR0tUjD0QW+cPdvTRmyIas3KAQ+kJFXgaqC+T
2qmqdrfysA+TXXQy1vxfl6QFXfLlDhP+g0+G55kPThjQs+iRrYE7He4H8xdq+uv73DCH/gZrBwE+
YRgepVl5ZuNNZbs6lVHs5Q/JxxMLoUejxZKbVsrkHbAR2AHF8olhjVSpXlttDEjmFZD1aBYQ6rtZ
0V+95cvT9uR1G1ZXocBOSW78QxkdE54sVH9kMLxPj9OEk0X0CTOJvfX0INR3CyJp/9Qln+nK5gVM
GvlR7Wdd8IvWfg9l6jRvwwrJBFUpP/iBKpBj/v4tlGHQb4mz0UT4Cw275kYNn+jOljH/TIfaraWH
pr3f3R9B2WVwNH5ZxTMRIwBsAIjvlNB1u79fcesbRGvqrX4KuoG11sqYtjO9DoUyPyspKBr8inQZ
AaE9wEM1HKuMrHprxk0V2mjfIq8kNKxyXvG5RDUBHJGFP4lRfCJExUlgubx+9gscN3jZbKp53EJn
iT0vMF8tHTcGeVjVnHYJW6gPAzLtzWErr6d/G/NYKk/WR5+msVobKRLoU4T0rKzNYT8gVqrXW6TY
BXzPAZTwNkKx5+fDVDPtFABFxkc45oUOdGlnTNOxJow3eE+i2+gwlpnIdGm8hBg4gQHrr+awgwi4
uqI9MWpcpX3k+/qra0rJGHUfBX6WwkwWb1Lldj8T4MPEN5L0SmHyN04ZfPAX0bXQXVdDYPhWKLXo
4pWhjCF+9cOqgXnRxOgaTrtqsr9Z9r5kTWBo+O2bdmQANByDguj7b8cPlwV0UXIWpWFdEF4NaKdl
Div8zQT7qtDWWIlUXkIxblJgWOAsb02kIicFaIVPIFi+afJfeFS+B1NVBFhJOv05eTTgOBR7P9VM
eP1mnyi4QPWyQLYjbIXAWRPeoMf7bApqyD3EjG+eumjGXx3BGr3eJJgyb6XKJS1tJ+3JXt2gcvDe
dtVlKXqXShXuNGPFQIswY4BHcZAaQIVCyGa+B2sGpiBAEXfU2OvnM32CC7CL1Bs6G4vggbfecE4M
seN2Ptv7loOu0KRegb2Mm1RZIWIq7W8arXqzPQz3wYyHoNmTTLnkMQMNr0R82rideav0vyAjKh34
2azGnDtL+QikWqLe7IMu1YftMS8rVfgR3q07xojNWjtkLpvaW7/Z8kSgvbIPS0C69VKO05VkBNdw
XFxSPyaEhux19pcucTbqNcD5xa2RoEIpVejsJMKpeFk/kb4i1P+V6P3a1SGlbQzxLNpZTXteDu4h
cBjRf9Q1qgy++TlLQEe9V3pwqC1IN1IOSVCCsQ/upoMcq1k9zeFIw7bo3ZOzfdrOPDF01P3xclex
JbLA9ixz2wpVPJn4fTOjYP7IOweXJmWvwFHO9OiEGUK+tq/mpYtCjXvHqg6pQoSlz84UgyOr+ySy
gYi1evOqH1YXaLEEpCLwJ/d4MY/+NpLYZf7wHTPaDxJhd4HPuIDGyzPct0/GH19tklRAbjhsCm06
l0Q/u92v0ZwabFOk0f011pbmThDy4MbP43xD2j4e6LQvoZsdCWajIHt/0X4F6sbDn32E2l57r5wz
bI66YOjdiLXZYGITMFZzcxeqf+j9bcjCPoEgvT6LSUzFZfI0eEF4oVYFU1bUA2//LU4PyYNmQV9P
g4/Gr12z7KTgPaQUwNjmGJZAnDbWICsozME3ELn0nzMkPl/vbDx7Xqpwx7rRo6cfgyKs5YhAI/8o
ajX6LJXBIX8SiU62sMyWaGbiOlztzY2XBNTxXoiodUXLeXjWA9g2n/HA1GZXz1gbZFKA2p5zfDVy
oPkuh/evNshkVcMnMXJbQmTbKWKyIDnu1IblDowfeEUsBNlM9e2LvUP6+84/Px0LK690ii3S/BCk
y6gnY2JlfZMflwL//v19rhNKp23x+3ahwizd69zgqFGeFg9GjAHsg9M5LW1TWxjsb5nxqcQ9rAzL
CC8zq1uVjugeM+tIdSilT1Pu/MXEEeWWU1NCeCTPb/v6GYvx7m8mniOdMBxoMpLqavbL8vKGFr+I
fxfm6fTBjErbKCKro0A1eMtrcV8/sn2q2Oe4dYfe7OxvhEmwkaCX4NjyzF3jR5IgR3TtYACahezw
Luk3ddq/VZ2KDBpzcdNNTBaqdNzUJM+Nek6NmT2ACX/Bc5CPSBB2To4sDDl52+ZKE7LecGXtcmiH
DD2NIbBJtwIEmtIwhePwDCcEcwNwwd309yCQeOnOMe3LMzYnpjhnZkcOeIALyoGi7Yn24DJ5wRst
j7PU3tqaXl4prjjuGYkKwmulX1OZMk7aamIt9N6IGg6OvcS8fz6RAfgN/n4QYUeRxb3tcSPKgjWi
1cSK+GXZMk4r2Z1z9snGGvmFJlIAxW2kFIXhvQkeQnjmsA4cwEx4KQRFwY5ePrFM1m0v+hhTR8ju
vIZ99/gWoUlLeFUWu7W8UDD6JmE89NhtL5DyrLe/SiFQi7p+k/I1M5ca3CwA0MQiblx0BbHdufBy
fYJD74dN1rz0X3IZjxKeK1UwkSi/C7qOlVVYNdBsQoH2vGAfY5WXW3cpopiOtBzm9Jo1VuwpMBfv
9lEONXttVoWxf7j9DvSIQYmxY5dKtAQh54N39KsJah9bqgmm19Sp3NfI6CpBlsuqZ6fhJI5a8k+O
JBP0xMgYeqUdoZm2vYtnrqTKo1G/3cnPKWGVrIAixCLXTHCiay3eV6/iKfJIb3JdFOz6JicNivx8
UfvgEwXMtmCQuCd/CgY6a0n2zKn1eHo5kpbjScZDo/VMb3oi/Ninrfou/fnspPiImUohLuvJsDSQ
ROr9Hh2twH8Gzl5ZNjw8SaDhMNmk+88cTlzm/gbrqWsRWLsTIBrlYzvOSUsAXocxKkUsVGjc/Ooc
FiM5qE305FB3O5DuwPNblWx6Ndn/v8iEB96bgNl9+waSGX9KCG8ntkjNjJvfIxOt44lqwcz367fm
JjQIvbuJh/jbCjeDbY8IV/eJ1XgGSopNL3i9fzds4T3CSZ/XVMGonhCDKtA80mueRGBZfdz+sY2E
lwi1CDU9H2LAwjH/aRm7jHYXC2F0cU82TTNIYV/zTYnorT8gJLs/OjADGbuHnOFja3DXB/Td5VwZ
QPbvafRAobMfFLS8PviPPOdRT+fh9qKfLCFwr8Vi+jifJFRNcGReYfSScyKVOWcitBmCFoVrv5Bj
+bHOZALKXmJ1Ykgb2r/Z0qHFifHo5Kw5o6FKi1hHAKf15+SPVabniOsFwXvByR8x6D+mGezMRU72
jAWw9ThRGzUXjJLWGTbyK/WOaFFPaI3fvz2CbWKn+HKC5aIRRqf3viNx/owKPpGVD8eehFUh9Dgo
dZdNeuby49RzoF20xgdlSLUJkX7lxqOOA9odqDoMveCQBOTXFsOzbjbahxLuvwj8tuDYdsc51xQN
rbLqtX+IlYK5gMJETFJIWfGnuQCMshkWDSa3ZO1KZWZ2v1LDlwjd1xs1Wiy6QtRU1812sBGXuI3P
XwlrbTpXGTiVbX7+mBxhOMPsEj26X7iHs4EZhW65V9j8W9FgbmSjOQvveFCuVDIYRcoS0B+LqRX6
xz+Qih6kUtIqxLyjVsWPtin1pTMhPy+KnrJ84XxPWSlV2qx3exEmlbivBoYziSogQD3HjOFVwIo1
4l6p1mlcHwJQTYsqf3+WYhy3l38b2sY/lAkBaemY2BsrgFgViDK45AL1qnSDbYl7+64ktkcd+DiL
OWFgtBm+6KmnMeli2pMsHifWSMcWYmqXvDPnct4pn3WMJ130IQ/eAVBP5VCEo/Jn9pyAvM624lpJ
yD5lajgqRNy6RWVYUaHy/A4ErzzRxl0+5c+boTPRwPMyNDRHeLzVgbIwI+WMyvvm13PHs5XiwkHd
6VtarsL6HxTaherPQlAxNHvweTiFam0Go+ZSufyHnthhxOdlNJ2fT+F4eTGYNNcCAqwBGzH/aC1e
v9mnfN8PrjPoQeGBkAhWuDsv0M0sZ68mBr/yk66Up2RSE1HHjVtEWvzst83nGfa7AMkFJeN09o+L
wTmFmED6CIjtWNgEJYp/E38nGucdoW7V/sX+WhKejHH4l6kLaSmirBU3NRqF46mLmAr7T2mPLwMI
dAMfB1FQ7ZT98aU52V63woBxUBQrj4LDdNKHC0i0vh81LXV2pnEljLoRNnibLxds7IhQ1Bdrr1zu
FZo9BfnzGhai2TSSqA0EY6eTyWeKT1KHnggU7V1defSGpLNV9HtUH4AeNLHzFGvKzc74kmu9lNav
NDoT56UNUf4pL2qVksFqk2oZTviyN5eey/5DahZW30zOeqzxhDKqWbcCYfAcsGKUqhpPbqjGEvtT
Vf+CpFdCszMMmm8vRuBYnP1sOrfVlm2xsq91w5kuDBz8kcL/ZhBqkI+y71XFVN3JVUyXzbqJQlo9
n1KHz7MgcGZhbTxACjyBQhWMK4vvwIUtwbR4gybIO3sNdHb0OtPE2hKFr/kGwFzgs0E48mOCG4YZ
FhZ7Ycx18Y2LV0bkGxdTmXlbVFZS994bh8/uYLdkNYDxkq3aFgPR5msyjofV2FP13powzkaKQrB7
00wIwDN/mKZ7fZCzpDvFgsoLdPhkMUNhvEQOSlBfFt4ppZBAQCtnCOWlUjrEf3IN85uuAhGvVLT6
ytM6grV/+A7eNu+OuxbWlr/yCGbA2Rqqq+x+Yngp1/hYRXTCoPlpOmhYqKxxnQG0Zk296OZWlcAD
Cd0yoqVuTn3PMORgbo2/pBM0U8dxxQXPlVgAo7Du0lm8z35I2NhqeSHYrFck1uJwvgyDN5Skk1S2
tj1edPOM/UjLovvUyT8uj/WkRHgRYLbWtZMsxMoj7tvBFhCUPQyxLz9R3AHUuVzqQwgjU4RNEbD2
5NsFhUQFj5kldZUrm+hG1w3exRH3Ywsg3R8S6z/7OdEODLq1qE8UNVjzzMBsHL/wpnr2I7lDaRTc
NA/pKDq0vGMdQ0L3lRdndG0dA8Uz6KbWzwOLAcf/pMMBAQNoNwzPV37RFyJQp6cDTOqRSDPg0JS7
jqTIbraPT9rxfdcdn8xFSydXVaRUttt4xYJD6pKVGYppdm5dHj+Y0P3cmNePcfzh4dwfT6rFmPUK
E76aePItrJlzr22eAZrP2I6beJRmGT4a/9ZHsAsu8lzEGffmHHsRyHJDks+QfL9R7j5uIhKqZ2Op
+c2dFJIixDNuZr0jA1OCCYwC7c3agYtrhBn9+pxJx07yh9IFqkjLCUizKwhTi4bEw27uY0AOkp99
SoZPy3tUi5rBmdGwkqXPyVD2aRgwz2MdFeYoasKl2pgaBsDZQE8TS+v3RVG+vPGOpYnawA6Fp9y2
IUlpYur0RWn6Tiy3Ot7QddbJqx+8A1WUInd5g5LPkj3igiD0s8BLY6p/b9gd2O+/XJ+zLwMibLKG
ski42VWCMq2bYxpMpZE0Urp1Osxh1hJ4Mv8i441fXA+g2LiAKjtIMlRdkipIQN9UrcU4o97joODJ
U8iML2GV7aDuaVqL/3IJYaKeECUMFuy1ba8SyL93UnYko3gZrEUGAcTytdOrUUvchtVGHGOwpwqz
XlKyoOy2+OSBpussFYEIkRrnSwZAStMZmz2zLdokl7nSA2G+KDbev04SUWQ7wCrz7xlIewEdxu28
h95SkE/xLbInbss/0lYOW9WCuOOFEkraN03g68X0zMRv2kSO8j64mC9UhxJ2xOF19lksoEcmklvf
8bnsb02+Q3vOJdJkuR9lbAh8aDwWl0o0ZPr+Vb3J/MyKqrNF0Gj3Rf/J1GThMq9hYboKoi5M0erp
rz/vIukrC6xaWgrHztoecO9xT9Db74BQQXYkW3crRl8qGPFtEidVJc5QtFbq9PyrXFg3JiRewUgd
oXKHUS8laOH2OhJhTW6gxP3UlZXKy3uuAqfJXyIqSYy5lPmqyLm0ElfVMx7vKRx5T79CEoueYL2r
m63C+a+6uGeqLIUveGWCujagrf2uvPQYYLjd2Q7I2ri5C0DWDkT1hnPD2j4TP68ytrTPIW005oFH
LCWii1IdVF+hyS9fjBPD9pwx3OGdtII9p7ZXr7/RN0dNpNr/xFWKLBGgNqx9qnn4ufQrovOhePvh
dYm5lWoXS8MOBW2nOyZAQfq8OQRdONK2TzLY5mdSUZeukwiuKaSlggX0jIiO/2HGBQ4tbt7GZRjW
jcnmx9h3ebg9WG8QekT/OEMkR86d2VbNQfSanZWJpi29HLp1AkEkg1YwXbSPsaurj7d1tdeyuxtl
j8hgUGRPfV6v0zJNL5r8u11Qey758uwwWwGWZWzB5xm77Z0Xb2Y4IX+enX1IvdEi+D0TmD9VBqnO
LoL5KuNXRjSMRI66ByNYXt92X2oc5PKLoDjeAiP3yYOBVpKQBSJHxH6tfXJzh7X5nclt23PnF//2
TwVXdaYkBwojBf4n/9JClyGbscSOjtLamfrGTvX53K3Z7QlkH650wqEA7SdynRqxPy69PTRZ2DAh
UGyUFdycIdh8Y5Bb+45XwXTPXPPspvNUhjePAXiPGsk1gSNQQfYgbQ9ao7rIk3PFt3xDlIDZUxIv
H6gi3jIt7l4W3G/0Bny4qaKXbnX3xuexBmrRP4X+MMpoDIA/I29626hC6QJpH8maj8ozwKhA1EjB
Q6nPa5MHDkpgiPI/akV/+3EhWrBnMM9zc3r+d9UD49VffBhNaD9PNKNt42E8U2kOS3tWkhqBGBN1
7p2Yp20TEk5FLY3zykonoHexPdQIOxVmMXnqfHNYvw3tq+AgJaXc3+zq3Wi7p3vs5Hk/xZfJh7p9
DVu7qzoG8unCRAU5QxBEg/d3bcVBLI+JJ650/9nIYvXM/P0M0ry0OcoEv7UQFEq9d7wySFoE5SVE
Y3z7GTNcellfxvtAuxrLybPOxPzznXSOVkCgjm6o1tJ1F7X5e8c+waGbstMfIeGBckIizWHEJRXw
zCRyUOX6azJS+XV/TGAZAAsFFuyPld6pXr3TKcCa8lt+3mc2qGhMttNEjP8rbdXHbnxBV9C9RmHN
Qx2i8gQB4i+zuPWq37kUFBoeceqYbH51CfrRpzssQ2cacptqAMp12Ijjv/Lpvkb7B8UlAHZ0sFb7
72H9qTH81IeermzdEUx8TdOCHroGsIOx5bFuCHZBA221jMfGGDQ7lgXRWFt/wjuqU4AqjH+H8WMq
jl1du71QvWgzkiMRzhqXgUADYsUxz9pGHJpUyO7RN4A5E+XCdASIobQ7a0xWZWXcfloYCKHUWIk7
ix8PoQOP9v05QSkCRZI+JW0ks5F4A1MunRTkvRMiVyGAMYrFeVnPVIRsFE66WdtRTREwZvKWK3/H
czPHFBwWfM0sA8Um3OhaMk5NQX8E8HcFXIB0xaDBFZ8FX7hIRfqfryLt3xDua2EUqN9w0GdS7NcU
7MYEHVH/u3PaHdV+8bHTSyRIiQfMwGtNYB2oorzy6iJlSnkcR2URyvVUC2Yq+tkUnmmS0lsuHJ7D
sZO6GrQBlIoA/th6pMiivU3rfP/2M6vuien3uMJP0iz6N1bCOX9yPLbFWlCcphf41Xm3PR+lwlMM
hyXRQ/+z+Vc9E45DpeefYoMOeNNVneZIo4DwQkHDdGhKLcfH3xKIqpw2eTSXQkLQ6m92raNra5+S
1WZAsxbweI4A4XdldsskaqaXMkODvx+GYmSHyvFYFrkylvG9fC1omS4UbZ+aYFBZuIABwfRTt4Bg
p48udz7ZPkfUWKc5lCH22BEuj6BfBRuLkyzcun+MFnnNr5LMdub/nmJkKAPQRlMdm/H4So5ttpxb
8r1FQBXptdjJTll7iTehLYB6UEjrNv+ZbGz7QrFMpIM7X7DOP8VWklUE8AetqyZWaVT/Rr+c7aAp
TaXpv5UhvzqnFju08EjTyKYKEeMefxtJ/r52gFu+4anzy9lj4x8d+0tGWXk3mKemIvgCyy6e3xmh
VLA6xMLO3lOpd4KNcpzRG2Rl9BEEYTYqV3JC2nGwhd6woLRFzf0y/8G9WWBqSmrC0qwcf4MLVc7o
jfhjS1IwivmI/GeYz7okWH5M07j356QpIJk2REw47pFcmuyH8TDKotCbcwQ6td5BTyntcd5oOeZZ
HAE0ODy66h/A7fZ1WTF+kRGpagCHlkTzb75TrswoDGUq30e9JnneHlHhWOcd1rLBn8dFi71O6s9b
OAsskhWE3aK7P5RzU1uaeViT9IeANvk//c+apulG61gBZtwshJIpvF+KhJgYYFi1ES7HZawu3WtK
IXFnNfbF1wh7joGYMHd7cr974W7KLlMiHdHdNmhAxiLYO35TyIvfjoeIRUArDf6JV0UrRJ8TXqMB
uKJgDvBZ9j2WQbB41CHyXmDb1uggZGMl8ZOPIDfSUPy+3ekddb+A9OM3i3DQw6WXz8zn6RqX0RzQ
30DdMZ0tlsLoK9+rNnrQjtoXk/W3XuLIw110q2NMvUu5l9ubrWDwqGEggG8al24wFsglPp8fhnmy
OkwViFnIzEEYr7OB7p8bjAtg8VKpP0B2Bmn2q0WhjB+sYPrRch78LZuGmA5v6BzSXEd5R6IRxTaI
aAvzgpzjo9+8NPRoRVZ40zFMeXVENHZtGf6u82aquPP+AYyYJbNN0B+SkAKiOFZ4mqg1w/yeoLZF
ByGz52ClaszuG0vMvvtTw7u37SNBF5yISq95HOOeeGnirq5P0Ehx8GEU3feHfC/Jry2MdP9ragkp
5qAsImhHagu6JS764qmMedzvJsBVDsep1O5uhXpFrH0vAwf51CIfkYoxEIYoDB419fZBH9ogNA0v
BrkdXJSSBWqRGaG/AcmvbwGEbrUzaKWQZHyt2EuS4JgggkxwaLfdNmgHkM6RFQlaYpt8M2Vn+1jS
uOYMA98uL91fSLgjbpZKK8XQvP9aaoQjvLt5L/JML8lDtrWWc603LNon2w0a5nfRWd8BMSVjlyur
jxvDpTYbYCxxQTch/VflbiUvftCsPO+LTHqk543qNGtZ06U/8qy2VZ3bBjx1dXvH2pM2SGjvIzLO
8brFQOXsClDrMfFDv241EGHWC72D78OVhSoF+1IPi4b55mt1bcsZQAXFo7wD9RnL/+1qAg724/+h
kvjgcEHXJOR1p0LTVwPpf2GDOpbOPyXjw3glbtddrmuY9Hi3SPED09j1K71vgFcu908WQMBOtrU1
q2aiDpHsfMWUkYws1ecc/ozdiHPyiXMry5fP4biYh5isb8tS5bhJcejnIDMHRO8mjuBG6jJTSF5P
JLjJPNhwhqas1Qij7XaJ+40NSYSp1/ZBSAKfR4hZTAX6Qv92uwoWuLODg1uhIvidCcEQ3KnvIagT
o2JlCfDDo16JD4Q5VQ8dgokVXvQLfA+M4ZMJj9I08xVo65MGITp9t1GX3PfR7bQE1xZ2yrbfIU6w
/ltsEGZZKaYIgT7N7pFHH9s1dTQcbSTWPallvNdt+jpWHmNrY4BRa8Z5KNqhqCigLqHga1VuQtfz
Pksgc88VrwZK3IaSIg70/+fjhX0tUXKrkEkvgxBR9Vl8Xcz7F7k74H1elMOTbBdzF8Jw2JP5bML7
/KnFOVR5qpFjpEyADwpRHde/L6kqY1TQrPO91NvNn9X/2gJ3F0p2t71jFw1/Z5dpS92t2V+37Hdq
aVXIukx0lR7HQqcdMWuUahE7grBow4SbJc5ii6ytVUKGsD12ATLQ+jmomgGfoYhk7tByob4H90vR
qXyPtsVIQgQ2qV3V9lq5FnojLS/robCwfA2vIeWn+MTjzvMa0dYzBXha7soEJLIfli+7iCT01Uun
VqPSIwz4RYYGTeZV9Uwr8I2bM2PPD7afPivDZiwWHN/4cnRkMi8xAmHALZ6oVnj5R4vDFbhqhuc0
bw73Xs21U+3zvZBBT0cp0FjbQLwuGU20/0TP3p32Lmn023OOWs8f2Mqhq1hgGbpHWECv1yhuqJgF
2ZDTpFbd0yKPZlhJE3LJF3/igp8yvrytLCMlcZPPHEiLI9ljF40HUwSFid35J/ANyBZiLMAaZG6R
X1Fn7SNWBs0pnXZmBvnjlAG/SdbIJiu1hnZCuO8BML1WdbKBvSuF1w+ZHNS5rQY3gTFj7N8Jr9kf
2md6J9SpM23ABzux91KoLBsrGlkkaQ7xdkstPR8afMmkk0tqNguYQk+8OpC3XdLUlqE+LJAfkiky
FEzE+8mBEv3B2pXQGmLR6+icviPFCoCL8kwD/wakYQV7jqnvn+gvjuYWuz3f2cPG0acZHn+l16wV
xNkWmQaCMC3g+T9thEsoFYDYt9zXd4IztzE60ayiBqf+ucBvRHY/gm8H0lQUghKeMEPDSaz4/HxP
WJrsTIb1LiBgNugDCWy4zSeNOmXkffHOatbiD52ud4x3k385Wkf7WKcPYRu+cKmdE+iNjY4ugbd1
oydOgyYosbKpRI2w0lyNM6C/hB/V8IPEioKgnwiuhpUFRDcSztIal3vgu97gN5dYPysAjIH5eWNY
Bi3BBjFZhIOZKC4XfT+Bkim1edx5AYqCeCT5TujAWYt4hiDbm8LTYzBZRpGm01xcX2kmS9tOIZyw
mk5CqZEBstgPGqjZRsc2B1mCGvvxvbOFit6qWIlUjHL5tfQZTmgl7XpXImAmRxSGqHx/En8DaO7O
ccg0Fq1oaawnwI7xFQx46W3hbyYuiJ3RVROUe866iB/XPVsDQ7GhllfCQWBbZrNuvTkCMKJT+8lj
eAj30XxViR+Jy6HEPSxfy27tZNLUDzWlw7+IlCWEX0A8wEBt4Q9a79YImp+MQmTxE83hcrJRGG9/
Y5+HVWa/+2279N6AG45M+u+0MIJmCyvoTraQkE6iLNUj6UDFJqUiamqc8D808V0OZXQUupn39OEs
5lMkvOwkZdZ9OHJfaKL7yjooyRBe04BfnmJ6Fm7e5tYBBxM2NcK4tDY6RRN8vCi6ptk1dXZ2f90E
udTMXWngcBBjJu9/yoa+DF0HOhuQd7FZw6Mfeop1mT6tuH8ZYlnAqsnkFMKwTl8XfDaQPHtS6POF
FHb/w5bP0s1dtVmpCsF8YHzVOJC01SMLNYHThwZo+0h7rn/UG6U8n/N9XySDdT/A9hW4nfyRFMwe
jRet9bVTy3veCgis7jvtKdnJ7vnjnJnBCCIiZUYZRQbMGNPAhleWMzWretjAD1yaiyIAwW1eKNdd
1TG1jM/uy8r/+ls7zcy531NZfzrX9pLcYtrSPRheVhfb3IVK4ON+tb8/XjwG5GY9VLlxiVYloc0i
w4mYwasF5JlNtuYW+l1v4emJ48KnG7fWBLLSJlNAAKPhUbanc4iMZgNjFiRk7Eyv5rS/sqHtqGAM
bQEk9N+ZjYw2yBTLrrJNSlhdJkojIgPa6jKP+O5LDPogKYHRgNF41FT32K8z0Nk3BevLxebIHIdA
pH880eHHTIOYT+46n/3B8xBNhuvMCeLD0i3geQHqVNHPD24dRjNmJvQrM1PSBEVvroU7olFrweei
aMkglE18uHb41WUfm/HFzyVos7Z/+NK2j+lSK44qkaELMDZsJBsukt/4YG2ezR1JPXbZHbh0PdsX
AyjnICu3qcV1VlD7tFuBYhNVL6asMBjkrAIDAc7j2HPgrHjzpKPV26GfLhC+a1ANUJSR+o451Kxn
qRMFrtgIsNJx0sLaJ9+oTJESErioEzJzNedj/b6OPRycwyR8+6h2+9L8m5r3NCMzh6vvw8o3ocq5
NoXmSQ1cYl7tO0hu1L3HypnCsZv73qbm7Ve4xWCe7LDpOrDgcx2LKqQdD4RXuVnwyYEY2DfhQDdC
M0SJkCBxR0MwYIAx2T2bC54w8wJHehSLwx06VHwLpJKfCneI/wFLiFnWKYEbfEzqHa5HhyEUlNPY
lv6blI1Jaed/t1DfYhMwEq57ga8mhsEpJ1u1JHNourbjMPk1fSmYnSOuEUybP3As+OJLuFDsszxH
WI+GSEmpqZs4EQGACK8DdIDQMjOonAOdKNIyOle1mQdgXE9SbWikIrm1zxCcyDRyA6TVzDr5HJP7
UCZJ15N8wcfewx6Q5SLedzmemvcD6nBN1HbP7N6sfpecZEyV4u4OqdMRcqqODpPZrjcN2PnWc46N
BILfdJoDjavzHFciYTPqjzynJanZ/HTVyiJprqLLCAFvtFGCGNIbiJlSJRaplDEHSioMJg7VPKdz
eH0NTMCqPgBVUrne+G118tbSi8/ZVZJUPpqjrg9UQbKHua5s3bzJG6wZaTRzQ8mHpMfAVjutgczw
Ts9ejG/G24E/LwsUjDlgZQOMHLy/W3VXGnvHGOsHOfPPzucbSh7fXMeHEoZZvpI6DZinZf4bGRfF
AXWGfPZWjZnhN5vRLtC9P8QjRRqjh2VgRRQvGrpbnG+qb23ykmeYOWGwNtdf0Xfh5b5stC3oXu1z
oOdbxvxzGTrvqygu8Zd2AMrjKqfZ5xpPpFETO/iF3pwqqGGiUH+M7eka3ijtvdJkrxcKObcNQjuD
dc9Znb1HfD6P3Hvdr4l8G3AUjUrLP3yBTGbCSHEg4bGO1Hk5JkmsJFVkvrCO5H5kSwbFcKjSUk/I
H8K1aPU6fbIrtFxV486HnrOTL/mH/ikVuVplgvSr3t6i9VfmDd2HuxcZSMgZ+hLtXC7KrcMJ6HLC
jrTosmgcdAPpKjZ/GPCg5HClBD1M7nCUBGRe+Ju1+oGYD7uqBThV9tdM5aKvz1CtHUc4ji+1HhmN
BZG0iSrM7VMUky9NaCotb0eLHFXOMcr1SojnRd+Kq89ZeAXdgalTVxGRqdw8dyAAxZUB6n6WQxAc
FDeP3z+MSP6+fsaGtsXhMYbk9fWOz3Y0dSK4KN+vkeCRBYoeem2PfCqiwQDK23eE/M8NtfpoNrEC
kqc4wrE2hGguY/UtMx9LMiiFJSjGWHaHkt+cpBbErUs29VNWYl6GLyFS/4ABT3402kFfkOukMtOO
a+sWBNdQLlg1OcCbIQNoAOuufbH7qyPgRZSf5jZVfE0ALFDw5zFFwo0nGH7pSLeXjq3aT2t4AoNO
BIIBvQdJ6RZRnDckjddB8u3mF/Pg02YD8ec/2w2AYNuMq5DQiyg12E30L214hGQj8wywBaW11BIN
MGmGtv5Mdd6IEecGLmDIB28co0DRMH18TT1X9ZVIV+rbgZo18Z0L/hVmN00rqczYyqM0AVXIWhck
YNrQbjoaXPVQwcqIeZ5bnjRjgTF8ZXjVKvajHNlo3tu5N+l/h+YJyLclZDTH7CVoVq3lL+gtePXC
sRhcikV6zhTinySPN65VSz3En9vhibpmF1hjOu2/obuHr/qQaCaeimmjgS20CcjGkG3GU/wSF+Lv
Kw6v9F0hAPNTHRGSzDP2JjJ2dVKPU8hV1UmATrQkgcqN0jrHNmJZX5KxFJPwQN7IzvcalR/e4zuM
9zVNlN/mfVanDePls0+A1V3NxFLCmM6ZOlni+VQL9CmslaAGzYmtT4lwL7pRZOuJhXL3i0uGOMIh
k3OUf4+WTG0hK9Tj6sGZfY3alUD8zCkvDL6qNUKwXdapInlf/6uZFtENF+4qGFflvTML8GqY7+7/
MmDK7ilNdErFE5VSZSWnRW3O+F9zeYqKblNd83SDWKdgNLaFTW/vAW7xrQpT742LbifMIKV3FPwK
SVB2YeviQH7x9+ae5vIK3wtFUfj7Hsdpi/fkcJl9WbpfWmMzTyLmI4zkuL9NPTW9LPpNaNgZf0jw
z6iure/qSE+BpmTAN0SYwaR/3fOk1v0n/M4mF1o3b2ZToNuNPL2BDvGXctz5Bj4UE7BZX2oFc/qY
0OkzFSNik3DqdPtMyCMAGYCGkUn3jdR7uw8vTGmauDFPcBYp9alQKUIz6mudb/Cs08T2dKFmhcBt
9tx6VDxCI+MfP6s1X1VNF6Df8u1anG52Xx0Sp7SFPrQUgeBFCXZ1DygL4Ep+B5k1Mh1WUhcR0rB8
PlckufStedaxXyoqtsIYmdUI2SDbIbtZZqbny56i816/vagcCp+8uCxi+4uj4VSXsvPqpEHstEjf
wuxiis1PCSgDX+S6G9wd3+5lYbY/kxnOBeOFMMReh5r2zp4ntxgp87XhAIvdve5OHp0DUJzYf99H
2qCg3MQhczmdnyiqyodheEIdaLUOMw3K5qPIsNaEF27/SPCVioTsToytJ6ZwO21tCiY+nbzC2GPV
LcUgyL7GJDCPXhjXQq1WjegwWHHx80qW1sTG4ivNgOZg5W+o+6r0ZUzrRwzXR/CxUG9RGjDtzo/J
tBKMURyqlQzGs6xCNt4OBgXMoaTwE0cy2FUg1dXe11ryXvqt1mfgukxsPdouf7an6Le57go6wir8
/UPdIe2qF6iIWnUfOPMbPMyOKr8E5C48rBwfGKZBNjnyauwSViyS+EIeZkHb5HkbbxvoK86uXP+4
JAIxcMUSksLVh6uuF4HMUznxyBWcn/hpY8KMits4JBFAYaV0I4S5XIAc2Z6AlMVWKYYnaeJ0kUR0
tM7da8JyTXZTVQCgdro5+Ic3wuool+AwrPUcTSQ7LixK3bSpKI3nNMBAj79f5PuOX1+Atj+zcQH5
4Qaf6G6ob7wqUWwpNOLBIYinD9s1xHVSoD2I5/hlm1VACZSdW0pTWPga/L1JVfQEX++hJ/bXZb2f
usxBijaf43cKbxeEXQwphSLlnwi9gpiLEcrbFJvpKwmO/tsYg2JZsgWVQCSXe0ZN6I0QptO7xqMg
fOYM1EvbttIaxmB8NkYjy0oU/Ar8KU93vk0pP0IHQLTlrqZNoT+ypusLN9rX6U7C3nNvfgmEVV6b
IjYjbKfEC0sjVtbJU0zX5nGACjYUaN51qwtHpnzHh6lHN4VWnYUI/DqzW6p/IbK8X0FGK425HwKA
CX3YC/figVsSVhrneLyEUF4sDYicJJD4zEQIHp/eE+a1OU3EeCfABucMRFQs9odZAqAv4VRnjJkA
sIiqSl1bszapnwRzgU/tVEHPCdcUWABkgyeUwij2VcjldQhTpCGvgtqaxPPNapZY+DoNPJwPwY2j
U/DvLG7xFbWjO4gh5q1flM+L/GC5NmdwUBI3bW+HE1Z0pryYb8HiuaWubop/Tbu+9PRhW0KGfVF9
z1/WWoSqL61/q1tbcUYbFzZkeK95UO0FrycK65D4gr8FDCrbSszbkD6KLrYWvNcfG5itiu9KMvK4
ShcxWdbET9xfagteaSp2/7lPymf75WQZZak6bZZFzCajXb+L0IXBHcxua5D7bo86ljDouVz8yeyo
Y9u4I+JT0UYZk5ExByus7uAvlyecm6lg7/rdc0Yl6KAqPF9KBxTcSbCGDgIxY+T28qO9Z1iU1IAr
MvGmz0fx9LpVW2tqjNv4tGOiZsDwSDyx9nJOmGleJ1t1wkVRRpmVRbTYi9LjIOBSqUW+31eFbcYc
iytNkaHmfnI7xrd1orS6ca60JckLOyAx7RedHLyVYiOz/slYlHZeb/x3tmJIcxW4CKdqSsSOrvAV
t7iZBH7u8zCqepBtV/arWLqpiPiU4Wu7VBvdUgM9NwMlmdSuvM5qFn7ABi3X8eymv/t1ecwGN01Y
Zff2/M+eRmloiqYcQkUjy6sZusWREm3Lr0FAIJuwT5j2Q9NMLtTjleRhtROAx1fGBS5Nm7WpTvg+
DHgmPpXgp+DMoCOG9jjySAuc62Nl8vL1vDERXjgcaLwJgqhBH8cuA6WXFtl1cMw9hWvPd6ra3vFP
s7RSGDJeQ3NCOxNm9Ll3lKIS2vVvFo1BGPh8bC4OeDtBdf+cGZN62pWmtAPgikhO0yzMw2+klsKF
AkoTMvWMlYtUucRMVGsMKOpAJKNqC5re7We5p7tVmJFwcKBAuYK0MWqnL1QH+Ovk3TVyTHrF7gis
CVPdSBRsZSkVAWjOVIJxdrnqidOqmQZr62g5Uz1NGVRHrwCY3gWIjIg3BPTvosL41RdQRwwtqZGH
dbNYCzVqclUOa4U2f6zdCs7YjvtZiPBMbuUjeMbzibaiZWJv8/bTSW70qzBGd3nqvOCDog5rfqzd
313n+7TV0k83AR/DBFnBHdZWJnY4itGuJ79LC6G8kVHaNvzqq1RgilVoWwvegoT2sVEEFF+z90xq
YSs367VG4T+aBi3Tn/W/lVK/TqkFcipwbgsICdlv+HV+5lQx45tlQotBn9mOnDJniIIr9ZiKoX8m
k9z9wOsDlzLQuVP9gqJc6zvz/2TTGGtoLP32Oug6SYyHVWViahSsKULLYYLmC/qMm3fD/F2AiHV9
BUIAAG1M2sWAkxtuKW9eWeC2pmQ0fDU/r8Jm85YVIEWhytllxNY8iAkxJOdvOvPBjjeQbk13mRQg
AkHYcXXPX42eE6Lk8zBcszGYGu18u2idVQaeWCMzrmISeE6VxxiXIBZgE2ETKUKHTmot0u6JTPkm
KoFHGo4BUmtKcbDtDojR7Hc8ssBy5yDRkafxic1k00kaUpZcEEArfPy2HGjrVv86R0ADVwiWSAzn
l5j8yx8YGWI90EaigVhlIWWr99Q6P7140ig2sroV/l3p+IQbrQwGdUqbCDqevKhgiHsxKj0CWVzb
uMI/Gythyo712+LslxvduTn2C1nuNlIx/tBOUCQ+3utZW/kwQuqhMQnw1FDOBb3FJL5ukM4FOEgg
JW8NQ3Eaf+23Udo+Tfxbtjr+PYMhD7i1QXVpLF5KReV9DQSO4zHZWGhQSf5mIeHdjGx+hHMj2Q5o
hVbLz69uAFV10G56oLP73ut9BHhDuG8PA5Bf3kodEEn9BDsN2GjuvFYh0bwh3iE3zTVCYDaE2jEv
WQw3AZiWYpZNX/YtDP9KQgzKAGb1WCAOF/0JAaOCcQfCCI05oXv8+Gq6M82fAGvF7JCjGWAogSDP
DbSIo/wWr5rxFRkTI0ImLD9m0rJW/WWMZhdODlK8hIIPieowScIP+V8lvEad/+LQ+i9pSQ9lySuA
V5J7Vi5FODz6Mj0Ea7rlcz0sq7eKgz66f6jhVmLqXIGhhu8d4Xn/az+P2mbu4tssCth8tnQmaUPY
1mADqB3c1i/klzxzA8Lhyl0VH5nMq674SWoJqodw3U3MkbIafAX6QrJsxB0iA+h9/qHkUckheSls
26d6fpUWb3jVeETeMOOP6GjkN1DToEA8UuchY9CRrCXMVSr31zSl/5LwMcIwJClw8gsW5sjSRyyF
zKotO76cFZu6gmEn+5pkyQWiVO3XIIvM2dUmacrPTA6+LeWO6GXXrEFtDRbxEX9UgJb11+ftOLAx
EfDQT8F5RM7a5Ts4d2FbcpA+O8Z3NvFxR1VJULSQHPDHoH0aGdO4/crOOmcfeVSOjXJ1HxDTKtU0
6MHVdJ1BZNuf/5Jmrb9cNmcCmM+i2Mtko1fa1DI50mj0KX2W3qHVwTesUuDnA4GLhsZczVQnPurQ
R59Vn2Z+ld4si4brRcdHdfRb2X2CM3c2mzERXxdclh3CeIZSY4qmwOhphhH/aczU/Bqz10Ed93kw
fd1RWlK+b+rlJnK56CcS+LSAyjMY51MI+6J5OBNUNgLhwCyM7Amc/Y79YcHdDNPAkPusn84z4ov/
7wWdK2H5Z3imtQU8dign/Y5JlxB7iC/YgkMzaMZBj9XSKXgXadaMzGD/gMaRkks3TOHE5wO+tuR1
Qy9six+IR2q8XortD8DwX4iMoG8wD1SSOj6wO+X7CDqAAFEDESx9Xl98pU/aZzDyEc+O3BwtTrKW
xgvyDbcMQfUwKOHhVAOfJ8DE/qNmtcFR6GjSHoVVsaLWqsLWRIHLVkElxyYGIkWg6LGvTEXt40ld
ijuWHbLQLUPDtawAsS4D9IF2d15LnxlBfgxggdkt/yKPPKdVKGgwP0bS2GLU3iJAOTzFbbVel6Q3
KQU021E5M3ooe/LsDww0gQ7TqPWBAu7GxdRWNAm0PyaNI1mnzWo3w4DhSrohPGKXSvsFVnJS+VwL
DwKDOa+LlDE5Ubbm3P2PnghWczxY7Y798auCqhzX9HfKUtFIzEZTR7ntXy3t3/FpiTCSUH+Grf0q
uVrGDaCSX1EFnjUeevnAQ80XZQLn/jsB2lqqgK3rYec8f4+bNs0L8Ps1YDJUXG18vhEl2thCE8xj
wJKR2ObxYMMHxzGpJMNEj5N8uNZGrgIEO2KVjXXmUuQW1edSSeiRNMh2uiQosuOvDiAESY9uRhQM
6iYXalf0nGTayFFWbFdoSThyZS35YUPyLqXTasVXclk42XEMTLJW6zq/ZGUcG1saXlL6OTKgMJ4T
/9SECBAlI9VrWY/xQTaUWlGT1DbdOI64aw4/KdIdI1FLS0X9d2fGoHYo1vatxTlFv+FtseRS283Q
t0Wvu1HiVV449u7Q0lQ+Lyk/x3dqYQgqzthpOYmtZ0hg5o8xF8ItyiuT+2isgVxD5RmaQMevssRz
AIU93uwQ8Wwsv6Zql45ldu/MOKpvSgf5ZY4YIxMqpfub+IMWD9bKKCunegHnaTkOWsntJxLqK515
pqIBRt/FakELLpx5/TOxXELOjAtTNCMDCM0Gpo6lD2jSMASKq/nFxopP5jgv1mXxyeuXyMpleWh5
CJeTgD1PwX6RaVjKGZ8bG4jGOHc+d79g5uV82UTcv8OVogikGfhDKSU9Qsvc2vwCTOggdWFswk4A
oXhVe3WHAPK3lxiX2N6yIrBuwkJ14FX78ywj1ss9LrO329UrKQjLit2LpD64UMJlhLtmihb6lh4X
a3NxpIlCxvDpSgAiiymy3sem4e2cbFmRU8dW7LpiCX6BKUZtrlOXrQn4VQ0kcYT/2z14BMxCJfYI
JmuciqsyjI72otZ13aYfICkhiu2Y44mTWgS0/76VnW7kUVqWmxRJxL8KmYUekCRHLFBtqLaHqv1i
+uyAoCdHdrxBJRT8GMCHGyIOmtKGHHfHaFeHp+nMFeFAi95ydLQzM/PopNa2sfmSPTWDhX8wrMIG
DSOaMBCciIFXCZHn2Is62VkFiPuaxjBtxRXjojD58Z4PuJVgP63eUOnhG7QfoPUrSSE9jY3AizDD
cmq7NFxErOp9rQnRx3U4utxoXGsBQ8Kpzqdy93iljFZ8HWEqEhcAMoHMdommgmYzKR+P5T9y0Whw
xxZnTh3K8QfvSt/KRwU9qIoB1nrTsG80922RZ7aWTR+HycQGosqv4o/5lZmyWBLcMGykRDenpUdv
VxBAA+ooTfZKQdCb1fd1tD6Q/LcGRlFLY776nbiiH5hVQ5xUWmTJBfXb8SXPI1Ox17ZcFffEhqxW
K0X/lkiwCSESroJ8iVNedqFUlHLpP45Thlh59p/GFIUA48h6ciYNhx0dorAgrsbq9yY8OkFc3l/Z
rI48ARv+ejlKTTsGz/fJQbwTvnpDanzGTsJsRy2DV7nRGeKoak/+k6adGLvOafEuzemEgd7jiJrh
YF8YOIYYB2OS7NXH4cSW0uel+QVE7XKW0fXESvG0rwaDfdB6vXXB8xhqpqymjwVF5RkBpOIaay1D
GHzFmLRWpH/WjLShXie58kwqsI9pRuZiZZwE+6IMqzDHsuey0cli/dksY0t84R06AiI5c//JvYO9
+hlfw63bv7q3YFp23w4D38WHazhVlAweJeUBcjEvFhfWxC2phZV9qQSN42MCM/xPc8G/ySNfvxjb
t3OmyIK2IECl5VPs09gAhR+dziHCPRYay51vHIM8CIrj+tRk0wIlXDbqnTdy3gbUPyfeaH3CgsSu
of1pkRSQvdbQzlByC0I7iPFNTH8+joGGJSgFW4TZ3xUrD+AUry7RX+D0X30jsPkCxqu/g/9yC/xt
1KCIluV40wrJqfDxTt1VXT93PqsBVMofrvIE2tJapgYs4Ll3dAUSMna0jpmneUh597CUMo8j5HYn
bK+oMuBLNnJCPiJQDZzd8S6WoHMLuzkAFFRURdocnysloDn2OxbAYq26fFw9EOhWnh6MjJUM3MHF
bjBt6uuOgX8j25XZjX6hWO7Slx8VEnq3g65X1jBVwHXWc1/bhxpYaOVWGKab4yQN3+Ei++Yq5mCz
y53GJxQazmthCtfQkzIqzSsF1Dgg46fSs+xGS0SBqfM3oTt7r87Wb0JieTFFLiTrZRWGHWwacrxp
na+oFmWpo2Q8CrPbfKNUfjWbVO+AEHlGitMu6sfyt7GECbYOYdfBqk5BU+diRH0Q4mlvkFp0zOW2
cb1hmept8OqG6o597RUBa15Es3eQto5DHAtdlxPS0pf4oH9M3SOSpwlSbBmcO76Gx8ZEez2r+JiA
RPr6YyJ4mLcjFQk1gXPMBYlqU7WdL8INnEoM994j3iFatPEnHaxhYqfI4O/j1K3yiHd9tJBtLfzG
BuV4yX7N/RmLtJJN9YEtrQQgeKZEsM7/YxzqB5y4L2gF51F9zUSZkZ9XuOUkkyQVceS/wZ8J3PBN
A6OmCaLIF9oi995MyvJ4nWWNIWip/q86mMYQtE4HIQyE5wCK4iJczm6xQqXYDQPTJxcn5cP+OV5r
s7Sc6J3YqpP3YQXnhaDBynwuQp0yDKlgQvlUOLPjc7zkQ6sFMMfeMFHQnkTBoOrHaFuaxxQ2d4NR
/pWHtYdbOrlq0Jz+kctto4OH38JZ+Qo8Y2VzAAMDbLkHgYX2CrPNso2dIw+HuLGqMgZhOJ6AsQxa
K8LefzaF4uhtmU8Zdhx2MNskqpLSPa0FisP+T5n62I7o/a4lN1erRL+tbPp8KfASwyWxDy2AUpag
Uh3ev4mNldA4GaL4cbyOLUzD89iwezp6Eix4EgjvLTtCQAVBH9jh+2Q8R0ea+mxAaZ+Sl9AneeFx
lDbHPxkUfAJ1rcOAQsan5NwlvzR/Y+A1h1hfT1ni0JL5IlKhWU+RRkAhUkgi3+oegYobF3DyEYf2
iM4PhWnUriz10McC2tlVoSlCm1DAYh6qRclZFgQmfiPR2kqaHs8aCXCU34mQKjIgy1phDR1E/v8c
LiceiKJ52H0a74qGvfV+hVFvk5Gfl5nyhygLQ7oBDu6EAkTWgEUReJrIyAzTvwkaqlWyxeKtwMll
si9uqOpzh7ZEwt8GL6ANRC4TFaslLXgi/NRdSzhytxKka0GlRguz6nkx5n2i3BFGtJWLPUJ9+WZT
W4Xd8HZf4pQ1oRqpwx9Lil7K0kI/ARGBtgHOrpp9gc3pk9ijXxNZlr7xAwJXxdftkjWEGx452e7G
gi1PIbq0FnyAsPJ52P9baOdL8HFNJ8PKMSX25YOsMp8SYYOd4eoFrQd5btx+rzzqYh6AM4M1Iu+M
P8h1efTBMmYu7jF/bSsSLo8lWqIKRXw2YlNpBPUlBpq8IVVipjn46gmh/tBcjjs24c3rssThS3HE
aVXBjrTE6pMZXIyNJ45hfG6jOIq6kZuXaAt08xjAl/v2eYROjooa40ylN3+irQk4ulb6Z2m/V7iA
wbFRKw33dDOe5kM4WN+Slr5MWo/zZbcP0ohVofO0h5COZ9jH+UqC8SdGubNhX+Z4OTLjXok4nFLL
8NiyDaCVFd3mItg0hFinZEzEBAzjCr12yIlzG6mtdmc+Sh9/Zax0TE7jXd5ZiWsuevYWsHbtP8hz
4ydKNVB3pikZTt5co7NGILG8GgcbFS5lM1kzIU5te/moKWhFemejOG4EcDPZLkXJjKDs7MQ6c7PZ
1vlP0NOGEcfMP69C9QZl2OrYxZHPWuCq0h5i4LK2sSv49lqD6uP7GagZpeKOk+y+zk9poZLuyxjM
rnE1jZqObpkmMbKJ9Sp/xW2Q6EyB5oPfMFWkC5vrq0z3BedhvLVnN/WF75LE7Go9y9A/6voAHTsw
wF4Ui7zcPwJxR6B8HFB3swYxs3lJd3JhRpFb0NbQKilipTyR/blwIY3JfKr44jtN5V/4cj8/012M
3tPOOW6nR/6dwYAKgp8xtwTj/Uo/BnOVBFHfMKWSO5RcThvRxZX6KzNGz4ZXptIMQyQz51UhfArN
evWRiqiY33FSALQBYyPY41SmltfWfyhMygEhHV5+y3ArcIs0ArhEfRM5egLt5M9IMfhTIUPi5njw
JU9Jl/BzefhoVydrpch+Yow/B2ElvIZk4zs5Let7c+EmrHhYC/TEtKJqpsG4mudww99Q93n9i3MS
W+q4RFGuwxJ6tTml9bGK7AfACtenqDhXRMGTqdquaeIQ+6E5M6C8jzR65O2NGTzyrJWxXnxqdLqP
1VahNlaKoiZCElSshjrNYvo8G9l0PQ6oJUtAdfim/DdMdYREe+0nyWddlAcAZ2yEv3VJP5/XQ59l
zlwcMYdG/gKkP4QELOG8c8ZUei0Ykpstnns3WJu8D2/J2SSfYY5i9vETVlftXSgoaeKhYsXOex3l
GWdkuFttyiH3M3dyNnW6b013uuqFBtKwcaYS4BxkTPo4mVFcwF8sXlFje5n7nwETrhV55RmMH1gN
/fqyZH3QSM+uJkAKwWACeeZGB8jAIBSTscjn4q+f/aWGT9dJtBkzkSImKgu7Xh12zQRIFwaMzHld
7IIpV96bT6rHNlKw1AW7GIJAOHzj03BtoqiZzgpf5OYGDYJHLVgm6KQqiPB7ZABPmK8MgRMvP8Ry
xGIXz2OmLdvoXrgAfJAkVbAZJaknf+9TEoO2Ke/Vb+dyldExcoBoADhLjDDV0wmfDaTOx1o5gMF+
9/PdwxsOYk+cJD6t8YhzoerNIEQt0bZ6zen4ywPLnPGXwr1aoy6CrBRCDmMboZrjNZ/Ai4Bux5Of
5DLCQWvfEf02LgeLnfTk4YY3gO12UpEAVGOC76Dn5zehN+q/qDUPKuiZvTwRfu8G8nB8xVFqEimG
PP8+luVjkTkY3CtvoJegd+vb9VxFm+ylJkvYv5VEE9pNiArZyTh05oXQmtR7PQCOkvxTVsd6CiEW
Ymg3TZ+/r9HjmfRFYl3N+VK8tBMfUw7u+wi10L4aETCfIY0v6TQFl79F+E1l+jEE62ejUTOe77zz
p2g9RvbuyFC5jBu9DRnU0erbC9RB3dsmKCv3xQmLJ2YvsTBhMtOfragVS7WNe9Atra6yTvrcQAs7
3VOVWewKAzyaOgY9hmXN4x1XwCbWG/YYueDse2CDFT8r6bnSBXp1KjcfDZ/f30X/iM2QxlTbIH7G
vd++xCgmn8rxOKZeu5WsRJ/1L6pl8QwqZF5mbLs8LtDlXLdMborHkqrI02VXs2cHYxsHbjKecLa5
Fiz4RXVVFfcEVVRsbyU2W9j0txxnlhk8f0kp9/dwu2otBmqW/iu+OAft1GiKEnl/iKQchzWZ0Oq+
opl1cUihT0eu5yehIpDcXcEEkRwxrMZhLPy0S4ykwPzA47q4XsCPUmDVPgWXBf3xYJt+xYI3TSct
n262RTEw2lWJXXOFZq+D4a++fSl1mSMg3kIJ79KcL6cd9rXi+L2uqW7pj0eY7me4lRMha8kbKLlo
sOFUZp270EumKpx5WZCQE0pRNn72ec95i5GvcwSN/dYNtUulXta4Bnpe2i5pGbZIXuTX/4dAleo4
shEMzIn7bgPakhXZ641qqs64qSE8WJha5zVDaO9xmPnRKmNZp8BUh5XphqGQ/bkrEBf5f/W+LcJV
kvpvk2dHtLt4TnOumVnuiVs0QGraaaJzyZLxf2tvD5i09bWKWM6fGGYzpt9tarMuHfDyqDk/aKWV
G9DvdJz6P1sgcfB0g3P3tZRY7/0GpGP5yX5+PeoNh58ILHxq8YhfG644WhpGNvZEyznaHt+2xYJa
HyxNs4lRLjcFYtO57uIQaVPAM4PdUkPsXy798AywbzsTzCWHHFjRrc8Rdi3xIhTfj6LsaeY8s4Q5
KTSX2U48ogxPc576hhqxnMRbR/etk+votZo2JhfSrP4fNEpiSdgs+37saTrC1Oq0a8jfnQ7BF6M3
WXY34DhAISo0+qj9booiDym/02ns7yT85dIb91BOt2BMI7d/h2/b5G29tvWCOXNinSFqUkFNb3Y4
JX+frXqljojN5eHwyXpeW9I7NOVvoSGZ31okG2dP6beyR13GprRKq1Y1NaLeX70v7OyGBrdrIgnX
k0A2oYWukcUTAbYFrOVim+PCL00MZfPCeWa7Q0FXDIwgMyukn73FEh8NLAtJzBBrI7G/3cHHGj10
zNKWThd75UX1EBHQsy7d9xTcgBCYBeKFsmnSjNErAabhLMAS207VtEoUMN+qRx2zWA3/VFAfoW6h
MtDiPWkZ6/tV7GprRlehBwFv3hUOGkOA29Y/ZYguiTwqbKrZncwfkPxkfNPNXA9I3eD+dQa3Hz/J
Kvdn+Z07mwQMHHgBv0jK5LUKeTKJQjEicAY16c1q/7Oe0gmDxvwUbegNRTrkbUEZuMUtLVQe6X4J
6KgiHfnq4X5OrrP1fkyFbtNk9LJhZ1XTJ9T0ywnAwTmx0ukwdZKDSu8VGSqgNZIJDCpF7h1qE8b7
lKUD8pjWcApqBh0TULUMOc6KhqBhaIdXzBaszP3+3ix78zcGkICtV8LrMYCLJsSoCarQNNkBsPSi
Krh1cDvftKVvcY7zzeye2zt/oJFDbftDTKJ4VtDfi5XlgsBvBQ7Hbg3ozJkAsa/g//h2iNCMbnR4
NjAcKZhdAIrrnYcJBPLs8PTb02nUF3g2JGtzOq3Pvf+g8ppm22DyNH5SOuYqQcij+xWMwczvvtE3
9jtDUs2lVYo6GLWfNa3FUxEh0a+Kx0t9kaJKKDrqsfFXyBIkftDT0yPUSqtPIn3qN0D4mGISBaIK
pJQQX0bfYpShVwfA3jmrDMRe2z1A5aVlehEqx2tp8gPiyv8tO6gEOHBfyF/u9e3xdQRj+CeBuh9f
Y19avkrikuEprZxTZPlm83/n4bOxD8nHzg5JcUiMefN5Rkt3/r7BhvwKyKRT25KtV5AsZHXCnF2y
p3OUkSBNxAzTu/n7E+FRbLE1OV8+tdpTZrCGWNJrOlrSxc/YC3aGiVT4R7Gl63gyVr18q5wljKbV
+MJzjTdq1i1CngpcUpchGCLCkt29GKY9O6GhL0uXx/u1opyV58VMhvTpEZnxaw6W/Mg6BWQTYLI5
0WUJhHzRsbS7trtNqMUiTDbNUtOHuoVzFYUseUvMkswx08a+yIQDx9AQusOzu84FfMK25c3zJDzW
hvjpf4zdnIbcEZLY1DA0PRaFHSH/bZ3qmSTf6EdfLGVQE+7kkXoLqMo0MBeqhkfccNc8N/pOxsY7
tybXWNl3fLej0h/qiqdDEft/DxXoTGbccuJAvI6LmY6W7tIzNojF1GQshYYQsqD/YDeACEF8vCyh
Vd6Wn6bzAJGLImrlla8dmmsJiXbepMBTtFpWWOgl8Ir+meZ7pTA5zuKX4VsaRww/+FkyDs/Oto9b
CD+ke7GyjvesNGga6iAUBbng4qTvR+rbm7tc6ROQU8dSv/G8/DLLBaIo6Zt/caYOE/BkBMTuaIO0
nw6PvkZ7kaCKtmxuWdF/GgHIIno4nlrz2ZryS4RZwiVy7OTlK1Io82DAII6DzHwDZch5S1ckZnfI
tYHLNJDwN1297cm3GUwZrwOL3cWb5eXgisXMlzl8dn/2FyIe/T1N3s8piW+J2FbaVORMDhMuC8Tc
lSg9Rn17Z8s72VDh0HIeO9mvphi3XBuYnPzb2xzgLgG1MSWu65basg66zN1faYSGxTTeLdQH0SBR
BjyLqazLGR7sv9Uyz5EiyyKPIx5G2hyXJnnGcSForwCrbCazFar68Lyxq+zVV/+AD392QBTGyEM3
Ak0zKuI9RGYgnoUSlv8JMGVPkuIt4jSoat02wyeOlVVbS24JgO2VhE0PrMV3xaB++WdIbKcNBvfz
P3ZsY5QQvKWmB0uuqbmHBxAhd+HTjkBW+cG/dIodVgJYzENYlmOWzxNJwStbOIddoQQgvYtR+Cob
WXCcfg3D56sPtKV0coxzXSsW2/nKGjbN80I0ZqlQz6uib7DApOdnexY7/toDNQOWhAOe2WZn4H3p
LyAPoMlSu3ovDbTcwGZdXIhgoGq1ktu7DCtn0jubUo9VaXn9ZB+7RMccxpv2Agrs2gwYZvmuPW5s
AK4B2FTX7vlaVlEk8FFK31Po2TIMSPK/nTssNB84N1h/3qnFMGpHRO/lwnI2mEa919BbCAB6OtkZ
BHnvkWvwvqgR7+3mJfVFFlXIPizS8suy155C7gNfcHJrbApCxG8ylpHg6+vpATMnuKsEn4qgkghB
Vo8sg123LukNRlocMaKleKhln1qZ4pACNN6uFUr5Sd4H2xhuBWz6HO4qMKF034wR/N1T8Xgf+nmu
PXGSU1EzurmZZ65c9yODgcAkGDF3b5YfkCV2wmUR42XGaczfclVhd0a85PVmb3wFo6oinGhFuuv7
wraGOpQmpqcIJ9xcTY6HdJmzgGWDX+fW897a31JSyWRT7EkvMClZME87T2uPxNI3eSpoowa8EDp7
/YUuvbTGUX2U5qExuUWCDjARcZI6asxplroXhUfnNdqHnJBgXfnkL6OxnNKA94xaLbEwnqYtjXyt
hG0L3T1xHqx9rYWF3mw/s2xmz5CRfKnmsLk6Vz4yBywInZJcpH+ta+ylYaejtxMUE6hSuQLi07kU
0DN0pxBuPcJXDSCUq9InB3Gy/ybda0lHaWtS+fJtJw4fkcbS/nFtE+aMu3QKm+iLSgQSlSKVu/kL
TQ3gK2JgA6FdXGeQTaacXzug7of7odki1LC+rkmkG+5d0DJxa/SZZ53BY2gCOgIsZf6W0VjFoF37
CTLcFHjgcuIw7h6OJkGJQ+Ig6ZzGuDEyJb1HYzXFnq1YmH9kUDnwK9ARiusf4sz9VS8m/d8Da1sU
Kjnzr1QHXYzJwRR0WbzS5Yd6NA3XqIptR1hDr5NtOtM/mGgbE+M3AaAbKgT4Of9POHTQIa7pluCo
vtZ8YFLdjel0yGaHxSDPHND7DfIMuCj0/ezXsIWfMCUYbxZDY003ku7qhnZetNsAsXyHti+WYKez
VC9QXHbjtaYJEjO9OT/Ow5bmtSl9zyFJkSs48zVxbjRRP9gmBHMEgmFwY/nVWgdOol8xPhMO3uoj
ybA5BZNGsgIAW3L8ufzOwhuQKbxgsxBfFUWfy5ri6Sxndgm1ya8BKoJtVcZpM6XEPS/4P9+yZFbC
38BQecmrAIn5T1zt5WnP/aTQEHKeivtTi1NM6vXvKQ9ZbtqnVber6nBYHi5VOL4MwqZrGqDwvrpm
cRI8lyhGPwG9BeCRBAP/iQC1biE0f7qURTMBnuxbI8gRmAHqQ0BtyIiR4rPxCPBOWAv0C0We79zz
yUKwh3allNn46bEyG4E1Wm8POxgF3TPb0PQVMl1zL6ySQpY2kNUTvHKRbmzJ1sTott8UpGvCVHiJ
EIqSfMy7CBTFqLJfMEyrgwi3gId6ixpQ8eyGd3w5kb6GO3ByMVWNG3VAnYyckau1TlcxPxxvANlb
imWjmG/xO44DygUy8tLW2YfLxGSW8MqPkyFmzbTT5USrRM8BUebD5dngdBjp2NposSQ7nGf3+Knk
ajfc9RBXA+pxZjJshMwDS4rauBfGOdcn6P3o+2nUte6z48FfMlj4KMTangk6IuWpoy28L2dBNkwW
VrMXjexlcFdlj9O5zYmsWkJp4IxL5KZbCqPbt6yxQXCANwAOgYxN14SgqpbeY2Pv+hlfkPji5QdG
BlFAh2G+uAHRPrXesxOp4B0rxC7e7FQQWoqhfpN6FW1WZuouS4aBjaMHC5Wz2QRMbBcIkPJt54PB
LI4Pdyu3M721morGluL0ofJ/4Vw+F5F1Z9ZVH0zZOCvVnUjV9sq9AZb9o3VqMsAGyyjJRyIG3BBR
xQocHl5KMVk591XvnqH5cZm+4p+YkhtPA7zaM6qWMzUM9X50lmCKI//dcAMraCkOoFxWWudnojrv
HvXlruRXpj68XF621NjkYUqoM5lpMpccjg9BzKeIb+BJBlHVmVBTMWisBGkOxcm/Dn65+jU/E2pi
YGcK1qDrUErYagXURM0eVNmqUtbl62XcuF/q3HxVQv77I8KXwJc0PZ67fJEkTZIpyKbQzvhzr0DO
MKqNs9+iNYBndZ8LigWwlRbZ/zHnVO0jQThACHtJXELEkQSJi2a6XTYUMmVPSQRIfq11tiYga+S1
dQMYGU7HlHBq5HLTmajeygF1KKg4PGo0IhHQJ4NWMhsbW47y3i0Fd3PW7zbuGzXk+irWo3CvTCS7
O8McEZ7ALgBIFEXoAmy+O+llPCgqTSsN1wuEGv9PEnhuhyzAO0hltCB51GbGltUoPm0Wdx9QjH2+
CC1KpAh0cPFS51nF/HyDVq70iXLwwJHXF9UjJFsqlh8VmO5tMJdP95oj5Ux4giSgOGIM9c9Aknz7
TgmWkIR97xM56onInxJNfx/IX5fpMdiE4/9/gRkBtTyHvDDMAuv6wE0hzPVCuSN9LDV5EBakdMNo
RYBJUUFjsS2fFblcoTR90W3XmD2qXXbuvocV2KQA7z7F0TYoOSCzM70aczyvK/lZh1wNxroknPW5
5e4cjsyVnvOOrc0BEFvETqtqEI9O/930ZKyvJ2Sc30N5GRdffvr4Z0WzZR3hBcgbwLhQo7Bffwok
Ma9y8fy6sMLhbANY7EWfZARfHj23f07GM58AfH6Yf/mY3fejwGA9Jz/F4mvV/oiQ6C+wFflvBUcE
KajZcILNj3oKHmRX83N9j20mL2BLKwQnjpkLy2jOcyjwb+aXawSO5jUT2fTlm4of+CjUumrw0J/4
5Hi4m3/LYili1/bQWtq9R3r913VkTKYLb5B5iu5+eTCGH+cRK+VIXxP7cTxHzK/Xu93q+QqBr8aV
XhPTz3LajraVyFe1criLu/peXlMJQC/Usw7dujjPMmVUAR95dac0D836WOoRpKbQuM2VMOZf1Jur
xNY4+OgFkLyvJe+v31b/93qD8oLsbxTn5B/3QGkIc1VmYUxYv64JK53z9Enftw6cYBmR7iGwJLQn
vFbCcTepxg6JgpRlZg5pkjkgvJh+2Nq8qxyA+Y1WKQMvFN76brsnG+Okf9SM4jH6GdqcksV1A7k4
RZUnVoMdNUKcvgIR5vwdkNWD65DCfxL6qJ6YfIFS6Zx+J7TKeD695TtU4dW0DmAwEnCAxo4NFHv0
RsRrBnEylzGGTCqOqCac9zK7f06OQG6DB1FORJ/3R7A9cTWiLT8oWBKTgVwspBXgeaYfg7ZtgeoT
LJ1hvSwe8OZSTwqq7El+7whSTdK6UgNl9dfTpc5Fk6wXHhpUqHK1/altjpt+Hre+AAKdzezNRls5
ZGPom6IA7jVRHa+KXxFRXLpl5MKV7AqqNRs8pQMC0tDccJsV4WZVESzOVRkruCbPpfuUbdQCD/kQ
7cS8ki0YszMOdFzGY3EFcE5JpEYuqR4o1PZVc9+c1dt3JYEDNbLBDExBE2uqWcHwFL/SZR7w+BJu
LP121SGUbjAH2rroliqv+Itmdnl/Jsxjh3uc3cY4ipoQb0jgGRLJ89kftu1e1uXMznZA0SlOm/US
Hqxb9wdZSQ4oYcZSW4TxRl3cZTbCPfsdEkWBTFYbX6Ajf8j6GVd4ck7OrEkgUFvgzCWo25pVMQLh
ZVB8Bu2aspfriI8ySRaMk4dfW3vrzFzApNv2hULb4ThMQP+HKignnJAfAcA96yjleCSRWxVcqjY4
kaQtM1tz1LyTRp5ejYK+OWAvj55QEu5PKtr/2Be5VapZdR2HUv4qOdz54EjFWkG9ha9s8Ea8S41G
4QEcE5O63ig90KyvqCsXUUtGHlNoemqEYTYnmzo1ZTjtfkp7x0q4m23qp6nnvR0/o7shPZ2zi0nN
vnV7jcPy3pfuPBvev+phFq5XOjrR0Iszzz2Gpx7JWSWvKDsBblgGa8PAW+Guf7lHO0q0BLaFMgz1
N9gy7QMouLG0g50G62Yo6YKRW2lMupab4T8EyEXf07MLSn3yf9nOx5TLQE7LYzoN/RSWGq6aWHjZ
WyF+ZQGDpFvKZeNoKhUMHlup4n9+Y90d28L6TiSPenSJF5T+/Gm2OCQqEW01T8plTGN7Y4nKgajl
cxUWHo71pseWNuCyp+8SIsbklEl2UniPe447BM9NsI9M22jMqc1SWDJwa3vD575yzMz1wNPyAryx
b+3DAEPEWhuq4I0EGAc7Msjhkzx4yo6ftwGpwZ4GNj2uGhZ4vucnok9rPfYdGfQk4JuzeVReJeMi
pD6petiKOqzRGele2LtbqSixfc2so2aEVPwmb0jLyc0IIMigQAw6zaBW/3cmq3bUhrCJfBS+GQd0
kzbHwThTJXlELA8Y1BM5xSgwg78VFWMWih7wXHqQsevlHIV3eBJMdHgH37NPwY4RaRrC0dHvmd79
/+CEd1jRCapuQ6ELQ1csTPFiL46wyjWmd8fEd/3W9TrLCBUjgVluA/qDE6Z5q2THLVjQSHf7KwMl
DOkaVfgs3IiRGiu79hnj2qzWD35lQOtd31PzEZ8XfwlOhg6jF3oaJ8B8IymUaa75CjKAm2BzmvHI
9CVNk86e81CbNMuOMbsVryFHc4SGANY+QIDcaN9D6nKqt+vkGYVOjVKpft84/vwLVJYxA0aSrCH2
wNs2ka8uv/lnNd/CxlLvf+uCh0xthfVGAGqDuR0wj2KIh9r9bHdnVXk5EED2ABhHJ/Sg5SCfNjrf
Zr9xvjFJSZKPvD5llshyIn9Ob48lGpCaORu2sqB0k25rVkpSj0h6kMRVVljMWH+m4+KQLuOINrRk
tc28nv/raEZ/YvxRo0UUcKGp3oDbv8PR6NXHVUBCd2WOVL/jd98EB81PNz6tFj4Zibn8T/RsIQ/h
I1QSjnhrOiJy1m1YxKyFlqCoVYIUtYLHqy4N8KAxSsZO/3ThVoiEDfQ3AdS3V4v2zb2caCp4yZ8R
JaIA1Y2aWQ2SvOU7vvwBdz8OO+xx6QyUxTMJazZoIJl8c1W5aOMIlJ8po4EFbSD4oGyie5T/vhcs
41VXewwWwsBS5z9BX6dNdtHtcPIfrhFJCiUviv3rhBhsaqP7KWjWmUnDMRrdtyt3b0HwuJob8IGD
R2IIGla3u24jjdkhqWNn80OequW7kHbCnzqqyBZGhu7KEtJLwL5z5cKd8SM1n3Jfrk97Eo7wIcSq
N/KZm6wwL1aego7gAGcONSsHFh/HUxqKAIQ+28NwWKjE2fX2ZoxPKSWNHJr8aLKqnw1B0VbRssFg
2VBVj1DUhWEOq7/LAGbdDVHo+1XRjn3spdMSk2U7Q8IfrcDRcteR2lEpLgNGmpjQHoTelqBrqnhw
JlvP8HF6PNdmdq2GdR21j85ZcYuXL+S0lrj6AuGujR3P4odaooreS9PYhGyS336SRtGZXUy/0+KL
fkB6Pty2I5+xU74rsvqgn7KajfnVqWIR5VyST6wDN2XI9ew03dcIhX+zWOdE1ZwZ2TK95hrcGI16
SOZTCWOrjrkzPme85ubnuokH63ZI7AdrRIwL5Qc4iQhs/oMP6A868PcwDVIEaWhtm7ZKHJbtW2KC
RkNSwhly4hyO779EVMBNnT1kUQBvv1INUgM585GQ0Ld01tCaM7hOy5vBke1Y/3JkUeM+93AmYSyB
tpoFyStS1GpfkTnmWQCElHdRx5EQ5g+y+ABtVewP0Tza1QFh2wCw90pN2QGAa5ZOOT0JAOrMvGah
O+ZUcjrazhUV7oBDM9QUPZd9m8OGOer0Rx2hl7Kx50wzm7ONXZpiztGgVoqyMwlebfCTql/lTx2s
mRiPRdY1yKUzLEFLQOg14kKHtUkCV2o4A46RphhlJJT1klyaOKSoAX4+NyrT7EfdXPWGLihVnHx2
Zd3Ea6pgr8jK70RpUDWKMcTuPoLlG4M3aCBKhsRTsF72dFu8/6y+MSPxSINZX73B7km2DUfi3X7W
enY7IGdZiwMvOgoEobTP6pYqYO62MnsuMx0IIlPdkLKTjNr+cv04FQWYqavPzUplRNarckZ/1p07
c6e+MCHJp6VxZ3Lw771E/bXHMTfwAgWPidt3VJDpS4epzPh6eL/W6EMf1o7D0UKNvGqxp5L4ZmPC
bnyISGhDdGpmHcyXnt9egb/B5tIxH3Lk9gCyIlgfFOh/fa286maYMZc/9OejcZVP6b4xVD/cpAcH
PxT1bw9V/3dz2wyg+PvluPWznQaFtmUNAezN+Sy83+zoHC1GQhzBudjwcSKEMOVn2F13EsWIPLhB
6WDH37MMzTcJLdOOgf4QyNaUCHN6PZsOeHsgPfmqylMQ9zC7Bh4hThzoKglEboUbvPJc1RrUeP7B
wbSunQtg7yQPaZ2j8w2wmI1bV9dmDVnFcLaOlF5GNKCTeODFyBArdzK+6/0vyP4KgXVCXBfesbnN
2576WqYQRnTi/acUXgeztG9EEvbtsDEo1Mbq8Z91lEN6i9h/7p2v2kv4XZSqZnnQ2IY9X/nKT6ZD
/9jtJ5tJ54bu8oC2azsi+amQbLSGFQgOJELye9bGl0X8xAihsEbPOlxmWLvUrPCy7r5gylWKUWbm
eTX4E/ySlY2YK4v+/Vt8cq9c/Wyfol6BcW7mwYp8x7pvn8AKrriRroWH/PgVDmP8NINOLQG1j980
gbzMnip4lSa9DTn0dXQqyXrJdmNzZm6nOFJlBvB5CbdI+66XwamjkJBPwja0dOoR6tz5KGsKdb/I
WCCWnnjx6O47F7eOtmwdblcGAqSrMJ1cPxh92z1dhDG8HmXt9Pg6Fm9SibDdS6Qm6ZgKA9opNzeJ
wMuAu+admqd66Hk05VKaqtXgjU3/qard8QMwKPNAmCq4gAAUnWhV7XuNDDR8VcpSmFo73fhf/05P
0IXIzD0WRYFnIuqhCXz2Ns557e0qlcykz3S9Cu1Ktg3Y+Lrd6j5qurtNu1DcRd2QNVnhqrrGAx2I
6+QdqjzV7VmrqgDss8DRZI6gspr+irFnDsFEeHV3NfmE+Fx5YTRGlTfIxTo/28EM+Fhcm5o3mhNB
vLD2yqtTO8GDKu1XRMnCimFeTpbRGavLNTk1NURlh0ddVwFKUeFmJ7xsxyPulSqw2RVeKnnv85Uy
pKHKxrO7CCX/FOaKZVOaXVWtyCw9FUqXqmqXisGrzPiJWI6ncySmY8MviWnYO1D8NJYsVrB8mdCP
44rR/t/qs9vPcLSl8frHN9OXBLa0v85VOcKddBc/fCLpcWssGeXFUImLt00KYB0XTicC16wXCkD8
cR+o+ItcW6ygeNbdzvuBZRscToogb5jnBAN7VS95BlGBDwe/qhcuSk6X7WhEYPvbMJcmv9YqTO1f
E6DdtGuZduZyJosTo6E6TeSdx8BQCcYnkiTQ7rG3AjBeIDBseYFdlFJUz7LZqc835XJSNXnJOMWW
xJWURqsnq3bYZ1HRF4Mjigku6kdctHPYIfZfLKGMbAgMUmvPEbnJAXhDyHB0JkxighO0g2do8uv0
YFu1uTPs4oxEHQVgbXJBO2W2ecfCVrO2TJLvYyIm8gtYLaYwCAkDYOaQJ3kv3oE/sS1sGvUz5B8b
tAQo9CBVlwacYGoWDjPYbc2LaY3ERpBT+4sFmb2WkC7D58ZgbVUaJmD1BgjxAcG/Mlt/vkEx8+iK
TheUhPGvg94Z+QEBq/TmN6RQtFMOMakG+oV6StmzwWNVqLgOAJq/YWZFagtTRLh64AdhzhSmOhOq
JEg2P7nMFYsNzSRklNmE7m7OH1RmFDZTuPLsgfp0hRb2t8lVC2xplyUcW7yaEBoowgmdW2ulpva6
pJRSdMzZ7c+IadmykRepYjxaxZ3K95faO1uRo0SASymXFnBmy+NH7phcSbUjnDoy3od9XOlOIsXT
4TcFNyFImjP3GCM295HjYkoux27zB5YIjvm8cPzuMyNnK3xABkbHgV6QlJ1P/D4c1CSpjeaAt9Oh
CXZOXgrfjYXngS4tASfErn0vhYKnoaKOmQ9bOeHVe/61JWvM5cWJxmoQ+QWLOoC9K93E8ng6LUtC
y2ZP9Lbp8NqSM53NI0Ypcgg2UEoTGB0DUvxPbkT17K4f85uKRbTZywhFTxlIg6ojLmf3kDl/Tvfq
kRtXEAxm80oAg6KLyy0R83XftihRFDVllCS1w9XiqvE8KcYfdDmAab8Llhbo3V2B6cgr9Sd44XMf
Gh5PxU9N+p1GpZ7vQfYbq+X/KNP1IGjUS9FniUjz7Tnei39iiY0oSdUoHQiisRC2fliTSA7ZEVc5
iuPVAmsY6n2J1yTkIOVTNdKgEPih930H0J8EXrVjAzGeKOyFabN62o2CPXVKa9/6JA1CkSpUFpD6
CMH+DddIwj3lx/bmgVLHfZ7ZsU/DFUicTq8UByfUFpE82PgpbYVXwIpxIkac3l0kFy5zavLClxys
mMQzBBfLYYZLwrUWfG+Vs/qQiHi0WaKxSkC/ZLA3xzrXTJP1/479hMGE3gYNTHn2c/vWuAaiNaT4
eDV3nTsaDujgPAu92oBtEnjuvbTcN2CWvif3tBITdaCY/RBPUxkl+le3oj0TXpln0mMSHc2RqauH
o7F51KSsUEO6LM8035vViKEeA3MMUEposufFXPstxQ25UYNROnShnxNLjYiouZCv3TAFmqMr4m9A
vTXjLR3HZUszP57Dr2HMVH8hKerH2aByQVzLd0k6KyNvZXXzVhZuvX4mwuIWCCe6Ck+MxZjznmrk
PEpMR6ht4r0oW3cK7Y2ZnpspkYki6h96XemxtOMnOKGki3XlKVc21sdGInBDWdG8KK20QrhIyeCU
DGOlu9QVg1udPJgXlEZ4hKJh51fUtH0MiyirqU9QJg/f2er6TVykrlQDOJqwir6f7BthtNBMNrSR
uxGV8U+nwpxbR/SetzSj7Ht9z5fAOEkO7BWyTIimMt3nYrAg6Go1l6JethZIOnsYFKT8WWHQZo4z
eYfDk5L4JPAb3F/OK5wrPDdd0HU/b+c9Yjiezr8CKQYf3v7QRblBhZLo0eiCYDXDwH3DuJfTuyc3
smzKFT5AHTFp6eXhxC5+lc6jZ5C1LS73SsJhuxzcUljSjfCujzYXQNGMVuzRneyopB3r48y3GvKb
E3344Gh1osadI+QI4IFr/oGzQbIsO574ees1eDadj8iW/nEaJGHH2OXlYTXhu9bfiFASsjSIs6h9
MRnmm7EhuIcZ+CTdboan66ucs47kwXNenrQ3Z8GE9GhiGAMGWLq1O8DCB12CW/yahWa0Q5INBM4X
qhZv2gM89+wJM4uX8Z0/QIUCq9LP5O9KysnGcte4WXqph+bD+T0XvQOOeiR0PIj4atfUWwDlVaC5
k9txVNAiLcQ/gr7uADvJP8+mH4ZC4yyPhVNR/Tmy2fnBai4DFiYERQN/AhHDpA/kL49bFeR2MrDO
Y64FDnz2hCRSUY9LUBpyDuW4+tbvRz/2avEWIGd1X+Olw0wHIdvbxC0l5/6veMvj4PgEyHvJtS5j
OzlSBw+np8kTpsP207tbxrLh0pBaGNCcqOsypgSi9HVMizi/qsaWkt4jiUBMqaCfEatCPvJzNXFQ
t8PIP8+n3m+tE1JvCXj8McoCJSKJr9VDS5/rOmIDNn2ssT0j90wEMZ/Dyoaz6Y1hJuP40k+JdR0T
isfQEinqNVvXCLao3NBLdHJafCXpC31H3BUdL9K41hF3j2leBh58ist2Pqa1opkvx4kspq+0r5gk
mNhtq6BwQw8e5bqhy5cGvrujknNTgx3Yg7FT3ibh4Lwc7qQ6DeBBHlIsSYBoTQJzKrMJ8Td3/9DG
Ex69PhcPCBkN4uaAb0m6tkqUNz5ruf2AI8DS7edbWb2g2utHFpYZ6EyJnc071X+Q1Wg9mooMBRSD
OhM5PzESet724PNyPcQ8aJAB49YCHFuJNaHnckhCjwf1EJsD1o+eU6zYsMr5Nqj4Z0pPoDWx7a6g
FKRyZ6uU6tmxyOuvd11LtkYxr6Z88Th2jhi3Cieple3B0k7DvZAcDFHhEfo7g7K0xkWp0NUsqJrM
qC4VrLp/vqI7h7ShMNhKFm2mzLFtPfGMjlef04qK9j7nCj0PWNYeFITEDKs2KeY4wsDDsB0NEc1Q
Tao9JB2NgUYCeUcSwFuiNoGqEIJb5Gm6D2dPTUZfQpftCa6x/FBnhSzybGMgpxs1wqz+Zu4MmheF
xPnBQ4YCdm3t8YK3ClkNc/wHcrYCFtJ5+vYf3pSR0vsUkWfS2woLkLq0WvvHlWtk0G9EOYzyGRuR
TJQMML1VunW+JoTVPOgVEedpY/PIDYN/YTmqEQG9rnmyAVE6i1pjwr9sFp3kNsVgMtPhtpMrbrEJ
FmFI9sjJR/wx3I6umeJcsc6yK3/G4y2VKeQoKoT9oyEtI2tj6F0uVLaFjAc1ZT+BniBQpg8nkxPy
8qMqbqthhWqN5dZvXpYXo3rTCmX+nIV9/3+m1cOo5WJad6iLOq9lA0LQfqi2sK/BQ6Cx2YmhN7HW
20sG+Xyx2qy+D9qLztWCCiAGazw2R1IGo7sHGhoyr+Uo7BlZAufdDlisJj3RGZE/5zjZ+f/07/gg
DFvSyn0GpTMt11cceNCMnGUXZzF8ssADWhB83lrbrd0QyMUC1ufVzvHOxK5uvU2Au7lLtOFzW0Cj
3EbuijdcRHUUAdqB5p1STg+KYuhEHF3afSFQHx6Kow1en+ab5cQJul0KqjU1KeSgwLRZdjt9j4nf
V9MGtZR2REoPR5ePO12W+4sAlu4HfQMjyO8GCwQPufpGsmSvbaIgrYQNfkeGAx4CTTv47Cj1XXmb
z57W/ltm/l+GOFdDukVptGMc7Tilphs/MmT8xPeu3ahCFATGtO3USGZIjgUZRcaixzxm3UtaphGJ
UJnv4h4HOfMGn2uaHp0GkTNQBRKYYLrMSWSnw8DgYUE6lRqAc7Icn0hQGZRp64pz/azvG1UzOxjR
sdL0sgnv+CYInsAmTlaHjDFkkeERdMT3lg954ixcObZ45GXaBjlSSntVbd7Ye143GzJY0Tnw1Zq5
AyjdEyDGS+GKKuQEEPfQkTzGwcPzyilv/0ZrH6DqqUR2c5fmaKQS91Il3a4y3IrLOZyLT6XrfhDe
vQCNnHSB7vWGqWayesHZrBxWJYJULM+L1QJSXmB9nyyaMr0SYAtAyJuCrZAhnuVdtbiWxYvQTW2g
xubVTx3RgYvz5aD5K27+sVSBOsIIrMTCitfO/FME1gxlwkvfV0wHCVrxnvHNp5FvJPHGnNz+c+E/
nUUagRHOklkMWBrg0q4EK8NKLjWJRA3i/n3BV3pXH8meKwm5LzniBcz+253kq444W9ZsjJjk9A/l
RZ4sXXMrGAsLqpaWVk97HnJGFCmK8Ii7XG4K1FILobU6Kgp/hkfcy4yMkBRFiCdiALQ3esP6TzNI
pZF14MSBYeXtDKPJx5omJj6/yDAiLuM3Ko7N/8UnWtw4d0gwOTl28HKz8xKal+aJZ+zUUjo306XP
olzvvVQqEnomqRHAsRS3JCTQTCXZo78OIPai7ce+UcnbBh8pIiPWAp5RYeRKbPaJyeh/WhNWwNKb
8yFIGjxIVSsDFPcWui0eV/3yEc8DbdMHfwtcTeRlbOO6Z5wpZ86g1VcyvoMGDWKOjnFPr4b0Xw3B
pZj0LlJihlOR8X6JGEe2TfuLEZlU1qETi7uU+aMvLw1GWhiMvfLTW2RotE7N+mySL3O85XrtqHhS
7hNhSXJR0XaGcCfhWdHVdzQxZXF1x3nDMVhO5OJ5vxnJp9gdKx4o21y2sd1pmkjMUxXzBVCWPyyf
TR6QGi7kbRKM5rlZGTl+ePBZ9/bko4mi7aCAKR7VmIW0UNCMyQhish6l28IpLqwg3ZW5iD1Y5Exm
hGg1Yw8M9AOd6dyylOI0AketdpqUHSLd4DyVWI4L2Xg5/emLvwEPk9UIz171JqqVBdn7tVaTmvb0
haj1kkkm8B315hL8lKdNSI3mU/Hx8SIZ9EyE3TOxv1cNcRvMKWt8DBEpjemy0cZ3LI9z4rC/8A4T
+ohNsgtGZC8HT5wVekLGJm/6sO+iw9ulHo1AtuszkIM2np0kx9d7M+80tE4TSB3bzygb/0iFAYRd
obhM+ZRzFBKqAqi+Rjd0E0ZjuLYHPiSucpErn10mzV3BxyGLalRH/al0OyZBM6o/J5YjcTRt8ioo
WN3InrcZhAnT6oKXjmFn2hxnXR7GV0Jt6WIKckq5MoByrxnb6IwTxqB+lqruP9tGNL5Iyv22Mt4o
yzw+3kblX8XpVjUAyC1uv7r5svhNl1CrPdBlCD66qFtybQAkQH+DlBXpf5nfaTBCAvndU9UpRuS9
RWwkWSlRt6TDhlN1C1rIaMAAqEfGpvSAEXJBYxbdFNRa0toGu4YSx9wlos5yloRfvwkhhoaJWs6E
Kwve9X30m0uRPbYAfLImwqW1ggbzjB82DuhkPQtbp0HtsQd/f1qGhPnmWc8VNqkZHO6Z6rxQtGN+
Xp34vkmW1HKApggnSR4Ib0U8uTZRAIYEgkv3RNjNsvZ+JvcH99qtMFQ3O9BjI87SAhVfW5R2utIw
MLuk+oyZtmbCGaMCnpooEQW5Xb00wp1xin8YohW1tWo+xCwVJ1s0DUjJdH1IEvmthfwCD1+IY8NP
D8ELhIn2SjgMxca53a5vkTAF1ps5pwm8y+Z8vzqW4rqJhz85jOK9JKCKWDep5H5LqHp/wf8rHQwu
Cj/FGEUMNZSmf1zSx1r8/XxKwIOrWkUO+fL2tVjBLwiZL5i64l0ovWr7QymwACOHxj7IyJRR3kZ+
2VnWj/7J9zVuBLDw7g6MGVGm8rpXa1rj0sVcuoqj5R/rFAsh33FgIy91CvZiM/aHGOq83CNlqeGH
VWP8be2QCpkLhaWx6deRXQm4NZdoFRROrYhVpEgBRlKp+7qn/kwmfxdpp13ZQLtmC0i5+4WI3BUE
xrnTh1lM2xVXr5JZt/nbJVkl7wNCly+odS9ikWG1Xw453gPjgMQnUQWl3wl+RF4qcAEI3GNB6RKf
4IVzYvn9J8oefvMqZiXYU65eH2JUI0DwjoDFEvADBGzIcdcKeq/7/+sfe0mccbpus2cjuOeccyvp
03HAZrO3xQxwIRqIv1QvpBLaBDjNOa4eMnAOUS9eEct1J3NWhs5JPyGCLDF5akVZCQgI77iVmCM0
KszcNlN8AWNxOd+Xw78P5TdidYnllO0HSlPplLb6VFJ94mutObpxSu5+CJwmjZDqX7vVfjT0vXrm
SuqfxJBDg/V+UyvB77RsLH1VzJCflLVhYi47AZPZFPZ7jguVFzwrCjgiT19IBgQnaq/aaMEpTG43
K09BymytjhOdT4/NbLnuU2UWzNPnaTjgOAjDnRlQ1COBJ4yK83veze89jBfzVxKFcVs8RoPx2uis
KyX1veyIQzY7uzd8GK+eogSXYK6F1o1vtQ+jPgOPH82xNemdVCwNPJoX3/AkfbAdqTj4WAB0e5R9
67zpDo4asjWeQZrGKbbU1HSfeNS3cSpa/7vca0wuBDS+EaAUPNkjTZe5oUan5WMjg8VJIYxo3C9j
YvvN1LG/q8d+EZKWo3V8abtLTfh0w0QB/T4QuQX+ME3cKECr2WpmJMjP9dU8DE3kfd40gBCr97jT
j9uI213Ym+B4QNHn6CscY+m75jhl1wSFMpykjAyLvkP6Xpy3he9BOJVkdL3youOIxQ1RgxMInOGM
BzcmPRq0IklfFcRvZMrGlruOV+mHosrcRNs5T+c2vSWq2Q9cTEzM0BVG104J7XT1bna1vtuSiWae
HyxpozFmDRHFxVdmYpncx7ovF/DiEgYV104rUKT+Kqcvmnmr7HpT72repDycWLDm1o9+JS1imLCP
B7Y3DrAy6fAPAynsNJUtnRkwdcEsycTzhmOYUpeEY7LFIkt+yJ5RxRJnlIzOPrcAGh5haTWF7Wz1
7iWikwNFdMsPkkzOh1DAPXOFd248rdeMBhHFynM64hF/PeytB+6GiOyVjY3WKCiNF5YFwLDUyhqE
0A4AT1SLzZe8mhGBJLQ1WApbfazCCEe/CH/ts/7noAfJgG24BUw9eRxIaFuVR6oZujK8DncArKHr
A2HfiSH1yzWiP+xpr8dKlGTho85ab4vtUI/asDbQoYJH4hC0vX6eV8VJmXdezhQiVWKB0mLyd81T
BwE112hFHyXFIQIpFYmXwaj/SVaqA0qHSjAUINhp4pM0+r9qDtAc9Pk8Tqk1IZOxWBxfsIfaUpI6
tVXHfqffg3FFdB8dmy6vyjE9f3r/PjudNcR4ywZ/jCoVh5THZzK4xptvaM3e7dlAAYVKbQXdJgiS
IHbmfkpYzg2jEuKmJXzJmIGTKAwGCVZWbcT2iCTlNcyLzO+LCQAehDmKpfv8Rsp8aWHboJ4dMt1z
CPsMYEutNhyL5PDKHr0VJ3hB6HBCGKoyWFT9IJM/yHsaF0D3KZm/YujvyXGpVlME6gAniSXNLzIG
Hm2iBthRlb9577aYt4bTqmMS60k2PCrqvcbjS1UJoPEC+M6RsVVZYtKQdizrhhV/3GXGsSd89CmF
u0qVwjf4/yU4eqqVTmcLsp2vs/RzsiLw3NGPF9NruvY4JX8xkzF46VmzX1Bf+1uVFvG5pV6fSgaO
k2glQ50f21n/N5NI31gW1OZAO0F26HBy2wNvuaIpP95lg0U/Hs4joRa70NqWfgZ1Ph8G1s4SpHJn
nDzCED7Pnz/gK/j2n56g1ZaEyQaXnE9BjahIA2tC33tHhk0t8EPW9jxAfcKbaG1/fKjDVUvRj5QZ
AQYpHkWBJkutDTdkXwrZTSEFNnmehHMuPh9EXj5Db0ywO9iLGOQ2dMfszieeLf0kITDMaH7I8zar
Ehk02z68eMmuO8q2G6fKKDgx2pmSgalG/ocD7MnQ9RcfExhaU6pyx0R1omi7hZxTRnAXO/ILWY1A
keALlZ2fx8Z2JJkvgKl+UDXypLkISl7793c10VDmAR3f4kXfISLneGTA1hwC/CkAhbvGZ1Byv7g1
oiyRT72JuEXcbY3jzJL1Y8H4+i231vaL4LpENoC2Ee2M0t8JPyMA96Lvy0iaGjmt+atL4u6LdQYO
RXA24HZe+uN1hNBkITFszdelBbYXcDJp9kI3vYEyLJoc763OzzdWpgkMvtpVI9hCUdc7yP+6k8Iv
O59cEtNQ3rUoBdzPAc7FJ//rn1Two8F+GF5lEHhkK3EtPa6M9/IDf0i74HiH0hJFqUfKLojbZwkk
XChkkBR1oEvD/5fx48P04BLx48pTSgQ9zYnBTy2yjQHAcNZ6Rk9uAArBBowzTXMXpZ47zm01huiL
2u8c2lav/hIQrsXem5A6SsmZmQWGV9rkba/OpA93FljC6/nsoPIma4FJ7C9pcrW7texVu8ZnDZ3r
qAOIrmK74R3jSQ0Gtt+3qn16mUvcHLs8V63arCBWkyeiZY1rsGuBmxcyuseNDpMuFMRtU99DRKD4
C2QMUiXIKYrSLu54N4YebxPBYZkXKcTFtJ7Cb+G8+aCKh/XPWbnZaOyXKEf8CLXZLsglAeIYVkOG
OYGzRao49s4qon1dcCBpXFop/q0qrY5M931RF85obzf1Xro5unedUjZz3gO8rIDlL1lIzhBPdBZ2
+VwzHZ+fXlPLU6+wjFzJbP589xI+4O3PBMMou0PG5odLIbayz939KOd/N3n1Psoe5pdkO0A4Chqa
X1CAbgKEh84vd8+k8/9Uty3X7lAX+fxr0xiHZEJ3cjn1dF070O6xzD8gxjRW0qNZ0fFP4fGAFKEl
YrmKJF8TKZJa2epX493N2f2GjqdrXb85wT4lHB+Si/qVJ0ps9dsXt6ZPrP73XJk9iaFaUF7+jHJ/
FsUvjGGcGvsRiBl5aLbzTV4KViterPrMUmSOoWUG+pf/wFCqYu9e6WlNIuOIQMHFU3x9n6Qk5Q8b
TINOQZ16xdOMFy/9N4ZoigF2WexrV01Yj2CDUJsc0hTlTkowOTpgOv48GpPElyZFnh1bO/dWLP4+
WWmmozqYnzjSo99IMEue3q87pX/TR7FaOooxgCE4hAx2I2s0693d8TaFwTIbXHiYez5Tkmk/rP1B
Ex6TwWZ7jenYziBBCT5zl46dBDUJnlUamrJB4CNyIIqxkgBi0Y1uwmoKC+DrwSymkt1dCnn0fWlf
cTAgOLJzMkeZfKtM47QKJFq2hzOYoh3JIjmWWnJh5AoQ7C46nYwqjp3nCKAkCaGdSyAHK+Yuhd1Y
aeEQOXr2yRCidx3/QgOzDlpvRzDbOhtTXd8jBQ1ECt9GymvtPM3j1FDjyy76N0PM3eQBNe8oI3Lz
rFu81H0TwxnxY7zIYYFGQNvKRYJRwCy4/5+qj/VLd8GI6YGNAjuQuiqrJAn29QY8AeQBieoISSgz
2iUbTN2NS3bA2FTlbmFxkEGGVAmreeEtuCjUmaaCdAtWiqHJd2lhwzJUxfiwlTYf/CZLdMGxrWYQ
+CpvkTCMrf7qb8Ba3sgWVFSS7G/ZEyV4QWN0F2WJ3eKgud7eciMZUoBh5gU/aRIfAnB6KIzK8ZHT
kgZAAyQxas6KSSxTFkv7WDKg0jn/a58pDHjvHCoFLvf2eRBsndqLCkLsBXfgPrACE0tPahlixFz5
AYY387thrK8McePtgb5gp0ey9Uh4Ebc2IitAv7YsPv9aRd6/QYFWHKQnhiSrYWDykj9sL5rfJpgf
3Wt65elLQk3yheaxQWQI030Xs0I+uW3LzO/jeo5A8WONxb6uHt2ORMwlISGg8aAUyd7yD9xkWuQ5
mRTcW7Ilreh0rS6x7n+Qd3X4T/qbTmgia9W5TKgBJ3Dg40SKU+knaYDlxXu3BNBT1MYs2sgamgly
vBc7NEzMkwnlrdVyYoasEX1bR85CKoOx0q+PfJRpOvtqs9arKZnHQqUN/mFsUV/b0pJOg4SOKpYK
DCbTwbAVEHhyoqgjejVIVs9gHf3HLPKWHB4JI/6hUgEx5Q4vH1VYE873IMk4R075/Dqwpgcv7B2Y
NeUyjJEGWlwAvymrP08+vgeTcu0/a+0SzLqnZA9pxR0oVX7Ul1VCJe80xas5T5ZiK0R2ENKfaJeM
mWit0OEjwtSVjAptrpAOhjurqsMO3TlB7Szhe7ZKXR1bvZpGjcCyYh/kvazUI80pW5SomIUNP/H2
ATWo1iWjvnskKavFMybht72032MfoC8vmXnO4w0iT4TbrHRaWJl6UAfJ23Q/Zn8/r1pirdrN5y6e
QzYIoUMnppDqHpUG8hpK3dgZrgBIfuUfAZU2tOO8t3gnYW9xXMjNV8ncU+ZVJKpwTJ8+5se61dlK
aET2Z1AV0+NuUIWFCCzzi69QCKGsZsJuiYr53I+JgeJZKWAWS7ttBRkKejwbIRJhDfPfzmKVissE
u7RjyNU9xAiBWSzpoB2W4T/OG+XQ2ob+Ybyc3xsJExC+XCihHnPeRIwU5Pe2Qk/lnQoqZBha9Xdh
ymazw4IOYakF+0nSPbXzN+i2j7F+dwP+2vlpmqaMj5XJbwBz9k6WJw7ItkipoZOeOK8+tABSfsTL
g6516FNIyipTFdq0vRM3JY7ettwgOJwR4VGqETvg3x0vqSB2/F3XWw8HN2NRXjmr7ku9KBlVxecg
1cWmqR6TAtnrE5+Z+gsz5etWoKjAMBf21HuZWP+v20A4bETrSyr3CYY9fgWaz50aeWMp96XIhaVH
DYK/MHhUJV30hBNBqGxfBenZ/U80xB1+S+9V7sBu+UjWSZR7Z6bZ3lmUg41+KDcbWd/bOt8gkQYj
i532/pqTdZK4RiGQ4XaXOEM3yYseOzzh5g4ygR255jFJwdDPrza3xC8I3yZ69ZyW6DkHDDU31PMH
fezwIYCHJrwVjMMpkzCGjCu4Hs50WX4vXb9GIEBaw5lGn1enUw8pmk5Vq+nqjURUJi/WEms22kLu
DmtWsox872LU6tj/pvvDnbW76pTqJIam3Z/dopwWFl+0P9ozLOJvDQJdklUxtoi/ebNkIEBJqQtv
j/6YqDYRqXJqiX0JEoGRPO7jqvxYOkDqWFLb5tlHYq2eTyIA9jd5axqEp/h5Jzc+8RDwFAjam/xZ
H5vTV06URyCa3l6qIp5NPs4HzdnTIRymCgqt1aXGJefyC1uyOheQimHWkkdhUATtXu628Zs3A/bt
6ZYmSK+2EBzUCdw+wBeMHbxk1Jl6103wsfHd03ExlHAdszK52C6AhSiB/g67Rx/BmRd0S7uRnGCs
aT/YEExcQzZzbsv4TVDlgxVqlHIgNvnYKhmDiFcpMuybFegS94571xaTBWv0StbcZJ/o0p4tktIT
l9urUFnOacoHFGP3ZP3kmE11hOhTs02MwbLlfzhCUtUQxFHxB5kHrhF3ahPuJBKas4aXGjK2GAAk
LpR3+pBjNTgYGN4eRG/wSTPlfNUED1PFgrgepUfJAksrRCgsDHXxsoaaU7ykkv35+ukbfHT82hcG
GRA6BzxaDFXNATp9U3igIPuUqC2luuWk6Cq9DDNguYpeRy9IiwIo+QniFcLeH1g+u1O5fkvSQT01
MyUo+zPOPVj8esluaosVuF26wFtWDaqsADV2CWQna24p+8lqGB1VHQPdZOr10KbHLTlQ8QKVyHjK
QE6LONhIJM7hwBC29LATAaLOetqv8aEE6rwMRjlpbi2hTbxy/U+2JIhEc3K73WNfKbClpHu+aIs0
6tgqWEFHjtcI+qFQEYh/yJLxXA6j1UnuQm/4pjlFJIJEsoC3PSvBJOuabw33hMVQ6nHyfkvYwMyd
VspIbFB2irRNiD3qrzgZr40PAcB4RzPOS0zJLz3ftw7fYU1eN/5g7W74h6c1rZRl3+0/MhhSSUh8
/xTbFT0b0uaNwFbwD8bd17XirPiiKz0U1sae+FplGuvCpVnlYfU7wQc2C4SjncZS6QitfhBCSjfa
IaOOt5X9HEXNTUVPkuLnlrdR9/xxz+BrJNyrB/LXXkNoovfXx4vlISFHTkuT3Tyg5TJ1F+aYaGIJ
rAc4ISkIZ32hV4BEFZgvAIqsxsXRoKBIP73hqNW9nyVWC+8pdxzdj79qbXq5K/RFKFHfbYSxL65z
nreUOR9e4TiDLp/7MrHpxxyDPblh9xmsYmWd8U5g7UAo+TFQoAIyeoUpsMrilAu0GjTDPPH34TmV
zGx2Wp8W2YA/l8kqr+5bNFcmKDFcil7ylNeAPqJYU8qEdVBNiwvM9dd1nVFYSnorzxbUF6HPgps6
aL6DZqjbAw1e90sS7bP4S6mOz7zBn1em77oD38Xw5MO0dg3s71wCxoxbVG+y93rfO0zoCWgta0NJ
DjjvRIlAELWG2sZlAf5zSP51aFgi8bC810tXRPCEhY4Ij1QHu8gfB13tVUVWrTDRcI1nWqMDNUZ8
uTi05oIKvcl9FYq5jDdyVGgFhBkAuKhHjgu1VjJkm+bcX8SXUAsIxjkj1NznTfRDdImF5tLxGy3G
pTGip05tL/dc6ohEtpxzSzh64FMF9hWQqHDvyc9LVxySTh/LjroISNDlMfinspBHrqYQLG6r+ZWR
AWQ2L2nTYQrndL0MXWQy9pYx6wuntlYeh7O+JbYCZHOc3bIyvg5A9lQlJUbkKGwURtCqDGs87kkw
rWP6Mdp2FGEg2LbB+WGFXnWDGDCLtMeNqWlucMgoc/lf9CEg7zM84SeDIeagj+oLpTo32VXMeojT
JbVHmbGBgnHawqtM15mFkOv76nSn6z7K64ipGz4XqcpIT1DRr+wSDNZ7KbBscvQJgu5pZeVpM5fq
Csz+PYPDPBSG8gwkqv2NZK7KlsdiLEph5GzZ9KWAb47KVCw8fjgvLWmgVFHE53TEEwgxvoMgRBYF
W9bkCJ8b2m6TOmDXzsX7j3VzoRcxKKWgQrsNvJK2yDSRALueuJlChOTYWX0I0RfBUaZdmsRkcwLE
RMSxeaV576qIjuKB5VRRzSeJm4H6waNFgFc9Qr85bYifjo7u3MO7XMf5KA7gPc5RTSLlSzNSjX4T
kkjYqRqsYYtAjD7uRxczkpUuLR2aUH/GIdyoqW8QJEOkckfnlba5AA4u1jT96mrafwm9vYEQVlaY
9O0n1CsFBq5hnYKxgaq1s6UFdUo852fL+NTvylZ5yTDB/sR2tOye4POXM4Wg7qm2dIdsJVtK168u
oTKV87dOwfAbZWqZUGCsbpNaF3YRMLSxJWxonCYRNz8TOqPVX7Exp0cIFId89CgeQ+yX1zgIfBQc
9p+HpRPZCoQkbJDgMqHN/x9Vhab3IRWKBsOMagEHNIZbnpNAO+9G3WoWpVHnY5IMODMpnT40ZTD7
VtSdkbLrnEBCKGqMEM9PdqHg74BZZNSPCu86FJN+a6khgF0nozzpic3pIoLXfQp4oMojx/iEqUd0
c2Cr1MI1zepXIDlJZ+qxoujLjbOBZGwwONYhmSv7Xi5EHk1ryu5No9q76OgyOjyRRSbxmbCBLpKp
TFifxu7spsB47XgLZxmBiIUtjHgMQOf1dskIlnqxn//TIZBddaD3R0I0LboHUGm/Rdnelr8zQIhS
liURrXThGUiHK9PA2KPK46kichm7kR8C3Nf2NLLNOHTPEdC2/QczSE6bhgkARDmGT2rQpi+hI7SB
kj2maq0kfJ+0YuVr/AYccij76mwbjBAZD0H9Hu4o8ClWmo1vVjj9WalP/09Omkn4CiEoRs1be40S
Vaj2V58xRqB5+a3PMaJ45AwEwtdpvXHLCEIe32cIT11Xbu3jMOc74fvnVyFNc4Ct7ZlX/Nv+j5B4
Dt99ljFFZYH1AJCXhmq7bz5LZGZx45slfB5pk9UFqEihVoWNP5fIZkL5an/A0a5kwWJPmBwVEE3z
d3LvcrgTaUBWzzX88eap5wTkP+bBYzzZi01RhIjXBNsh2hRn197L30D5577ZJeC2RyAK07CzJD40
RSdcPf5s1RNOyZTnvIrmZhfShdTQNqGAFCNH6Hvct7hr5Ppw2w5HCfJBdNNJtB8T066pDALuD6km
gBHRDXd+7S7NkCPRKF0Rir4SN8O4tETrdV8j/V6qPhpQ/pG7urEvtprktDzP/FChl8bOrX0RELKG
moPuLjs9WTOd5cX7lsgiaGVKI3ux0rnXoZ1/QxNaAS1K1L7HHaIRWsh71XJd8kKHCSCJWP5yMflk
duoyTP6RQSKZi9OBx8maz//F7rXGHIZ74zasb9KEvtk5dUNyL5QEHE8eHEG+CHHz0LV2Hx4VC4Qs
Bb4iL6AcQhDWxnW+eBNVITbEQhp2MQQgfdQ1xV8wGTDYuGwVz9vFG4Q2JLl5EWSc3BYF3jF4uOof
1dEjSeTNwgsN9RZmdCEGbRh0l9UQXbljxiRJQcmUhRIays7rzfF4zQQ1mimxGibyFqQ7glUX/ZxQ
LbjeW7ZelFMa3uY6FRlqf5g3NF+hvF3TIGQ+Lo7fvHOKGM2tu+jK2Zc2qHw20yY3i5cmFlRYbSkk
AOEU5iSfORyNkaKxcXVeSb10GnJnb7Ei+AMcRGBjFDDRkGcAAhPF/JkwcerYVHTRvdsQLnzZGXAo
mT9NmaHZoc2im3ZwMON8ia/OMJu/DzXjg9jMg03F7te9dY+CiSelXEjgEUNHzxaiKuIlQ1mXcWtd
yddervb/0W65w6LDDBTubvbxNhA5RoC93MAnsFy98GSV0tInQdWIRWi+lXOXUlJKyI88SxHYh7tY
1Lrl4Nzllue2HudndAN4VmE7X+xDmsmgjgpF4L8VxsUJs7n+TfPiqPubmy6QWh0eadJKL+ulGaeb
sIr4T91GbROF5AZcVOeJY8NBFuGuf0/WZmZH2tj4t7VOH0C620FrAFc23Qrur7mupdQ7euHIwV1o
9iSkTvU3FJmCKgouAj4FHV/wGpxKQ7v5PdIdK/oQ2zGJcOiN29poQbVxWXRRgxdtyrLO37xA+J7S
lU6zkmOpdQgUgW34F+FT3XDQxc1ZuWUtcrnKBt+oPsnSAd5gqYN6mRCl8Lka3MVj55ADe+ucZQdg
dpP9zABh/mWj+EAJ33gue/pAXo8ARJGUX7kAUOv8cWwqyYWDXvb1E8GMxYoxDXejRIGbzONuwzwZ
lTQ6cVy0oiQwt9cK0khdnIEohJEyxygsuPo+qu0swD2M7s8vTTNTJmuUbyGRi7QrxzcXZKvLaDED
Y9EjVbWyiBGZRoovE2W3MLOhYAbUWjefTtnqihU/FDe38nKPYWdjuFWq1KVCyE7rpFe5/oCUo/T7
Czl/nF5v/ibTvTStTnt45r0EQwKcQRRBTaJWoVsR+lYoWecCbvdvYt4pAaM0vpENLsRo5/dpwtCq
tK+PRxTsnRCD9++9rkcZvijIhHhj3BhZDzN2y3AfbceRQ29FvEnFwh0fhZjLEDPvWCoZAeM6Kmfr
+UOEBuBK6Cj1EoIDdVnFYRPyNFNkrDD+s7b+ZbMVV17Aw856lM35jc6MTlREZ4zX8IC/ZBj4C36+
VyCzZJjZt6iI5lI/3daoFxaIV5petFGY7q0Kna4J+0zGfcwLKDgHu8vA+KC1GiRFvRqkjkPabMo5
YYmAiV7mDvUwow06z/nI51V+1wXStHkBl3m3YiaaliY1PT3LOHoXd/D1QtQzyfFAACOtTGiCD3nU
AeokCDIyhtSk0MaxXVRGMkpS5pPEiSfgp6N/B2JiYl3RyfGBEYFMWQVH+W66+/1xyC/POadi5WaE
QdIc5FjyWZR3txZRWOJF4asKL2x4MPWKIxmOPG0tKW6yc4rUduiSEAvGQd+DMiWqfiIaFrz0Pcpr
JrnL8ThhRE7nfrPDFSIno8Go8ewTZIASp4uEtYuqLsq1F1MyZ0teKgUuBUvzFVCHx9eInVtpumOK
wQ8Xru31fNOh/E1XI4eCQrDuxqNMd5ZPVf1FAkp5sdOjpj7guAvFV6TIXFNxM/XLXUZL8bZSKEcZ
6AD8U/LuSNK1i/21lZBcIa9olcttc8ndsAggDhl+4zcGsQX1gPIa3eKRkTIyV4KIqSuM9jr3rbHG
oz1rttMhvRwW13N9g63IqjIdGA3K915r7aZSkRbIBKoX3CHRuHc8VIusS1dhWRTmY7BNWPhsW2G0
cJnh6jrzqlQOAjUM2baRp0h0sdFEd6z8ixXUxFiyXGo0pVk/ADqZjZp4i8KCdLyPzPxYrTLfLDX1
Np0svHJ3Z8k9YljmhX2l9XjH1xpyJDrxBDxKM4w2GStInMfZTniLlPZxUAVOBqfYIj/BJnLn0qEu
0IwjY0bVxKwMiQA2apPmGl+6yG0ScFl7uHS34bTEtRv19/D4K0r5L2ZuDZl09aE1mYLbsq0bU6eP
0hGqcNWj2WatEEHVn+BA94r/0iYI55tiZc8YHJGX/mw5ivFXdP/4xAPQ/rpiu/3AEaunRwCngvGu
Bt1qjKLPeAI+3DXlO8ctu4Mk9p5bAFtC0B4Zc4Gk8cC+UVb+7NsvhsRpoZ11gJuCtvR4tjCvyMz/
S1SGs895nXELW3ArZLjLpBFWDQcviVwTZCI/s4u0fApEW7FoHS2UHCvsH/Tr4KTbUGzSAxXypH2R
x+r27wc3aK0+JUUc4WnpcytP/w4r6l5k5HXEgahlkrUAnI/kphbO21HkhmyhRq6dMVWAo4/kPjmh
kemB3J9uidalDKT8C7qi/SDDKJvyzUQlLcQbmimD8oynP96GsspoyTUYCxpTJ2yDJNEVViwKxJyW
+l/pqV16ZH26KUiJlFpREUvho2mp9RaBZTlISsKzpuadvptjKK51TcpQxpw2sxfq1BxpF4G1KYL1
JBgFPsd1Bj2WZ3UbbJxcYDp2XS97ww1v5AxwEZIKO30bFw+pgNkOGxRApx/vK5zNzIbg2q3W0PUA
RCU6qfc6U113T9FiBl8cWoVe+/BLeIvHltelMAIo7iIbSAiZi/enGvNhruVAeSK4+pQili0JJbJ1
/IwWDPBKnnhvBmiRoYvu6Shd5HmHyuVLc47NYP7JNK8fLOl19/zfGsr9fOwgXYmGfPPUR6wo1r3F
kqNPZytbLsWeRcNibHkUkQsGYyf7NlYMQf+A37EvSmF2LRQg2ghjG3Twk/W3IZ/gQGw9SN2zmD6P
M+4EAv/40xDqgdbM+GKvo/T25nliqOQFlf6PDcN+DC8/tXiiql7zSoCv29qd8jomGsbLevIhqMDL
ISw1NwxhLTZK6EsXdOSYBYrPmOnn+Xg8Sd+rzjsN8MXeXIpCjioPGFCIezDNOPCSixIJk32XIo0q
MI/D/hz7pA0JaAxaoLkSxpdcKAWUkDn58vudS/0KqAwUpXLL14Tl1IyQnDbG5h1QYXGQXyDCsKq0
gayfzAWJMB62gcwYILnytT5wE63/P+hi6jnWE+41oify5EMG3uQUatOqSeCw23VpkAQsTkbs35CZ
qb7TJCPtnWoTBorZCclPqp9ECxi+X2FRiHPW7YI/JI3OkyY3MHJBa6jHhrpe7PhFwEWSp3Mu1NnQ
xjTcipO167RyaO3n1xvy5e6STfyTLa1jzl6xCbHTriok+Dl2I1nZ/PNAOWA0NW4qS+G+MG5x/OSz
SLiTzNAC/t9EV+iJ8z6JDnT5qIbkJ088AdYY3rkH7NabtG/3nvNWZrvEITXatzZzxZOPlmMEU2Xf
sJ6LOdN0zWcmvv5Q5JP5eNVkag+YmGTl6Voo4OOM4nJWMOy4/OSdNRPjHSt8XFQkRto44RRY5QbP
o9U7Spsat1h/Jzo3W+fYqrizv1HjToVgQL53WugBvSUmif8M099K5C3AUKhKQlz3UEwgPwTN6RtM
rORhYAawlabf3RRYPUFLFEP4JvN9gZZS4jnmi+KDpRJUDAG0BnPEYdSfDGj7PCCIePlNVHJy+oqT
PGvbNf7xv/qKQMTu9e1qhzLeC1uMJHYYFm2kbW+Nq+ZNlwx05AfHIoeQ27tDOW+hziLGG/4fTo2z
6t8tdx0q5dKQRGt5dHyWFFzysuWe2FUtWccaHa0xiIVpsBpqvH6io4MQRYBE3Ci5ddMFdtcnH15n
y+zhbmgJ8yo3a0D0neQLp3CVr0XLmFRyqywkrYCZEQGNaNX7zaFfH1QoGagVmPqWizw9NmOJG+8y
IoR1TKy+kw9YR6AvNL1GlLjc4xARfzo2JRn8vEB3OrUNgJDK7KFk6iWdnsd9ZXveR8zOjEujfxOg
wVsEnBNNlnNBleqeX/EwSvQ/SbG/iwRooZdMeeNYeBmpPjlO59i64upP2X7EwIIlaCrIZ9vQtnIv
YBu7QwLnhonHlWU+cX37oXlzT4WXysZ2xtJD6ZG3ZBqcYeVSwzZApb4K/NDncjh6jFbZwxbe/0Hx
sIf9MDVXcJgM0x99YFbplaEosQML4ruA53GMErL9sevshSXQdqyNie7w2esn+BtDmh1/pN41u+34
iIaK3JF/IQ9hX8BMtEnkgXugtq0pgMIOovFVdBFe0jwDB+t+pyOTggIA/ZRdzdPjmEBhqpyg+7up
gveQ8wGdDCML/MZIqUjbKAIuLCU0D1bVnI8vOyOJmfGjnFnfSCo1rgtkNcOR+4qTp1Fi/e5BJ0Yf
ceQj54GTgGb8vS46oFoe9IjoroBz9I9iqiXo+scp4ZcatHDo4LuZNsS9gQjriF3lzo9a97jRlUAL
ImEE9BeDSDARkTnFXh92k1y68LIH692LuGcPmJzkwjFqJ1Lhj+lgNThqLKSw1uAy2I2nY7/sP1Fx
BuFOlSRrKQrm7kBi7w+B4slV3qLizXM5K+GaTM2QveqUfxfMuQ0oF4dVjpE757gabYZaz8lZmIf7
kRfxFmFfAD5ETOjVZcvR9QOIbxHmX1Dk3XoessRoZP8LqsHaA0BfRozr+8nfp1IbE8f6eVil23/X
YceoMbsIpb1dwG8sLRB3/+WxJfbT1EVaM7r9v6BKb5WGdt3eJsCBRQn/lc3U4aWymU94q+XQgO2B
cRtBLxa2v2JozupOXWYjVB3E3UqA+OiuaV3Jq/A518m6gIuOTK0/aDUZO5uo/QVRI7QsqyrrvXiH
d7tS9JMNj1wYKJDOGTzIOVZKi//gl0CONE6tTY2GUCP9iQGrWXq5t6GvMKrLh6hkT3rIuxo6HjSV
B4BsG2e3DsTawBUYYnuHjqY4hxs0zAEoCpez1viEdyh6i+QJqw/vahr9dODgw2XDhh5Kde0XznU0
RWm/vSyXdca7yJEWbfHu8ycM/JzHY3mOFE/K/9H3AYEas9054fqhwgQ5MwkNE+mUQUs2bEMIUriQ
gZLjkwJG5K3iEocL/SSH8pYWx4Vcf7WtorcdZVPHWPbHz6MxodI8P9lrwaBHVTs0e3ZCC4fiVlsC
WSWd3SY+G5IRfNUnQOT6k+clfgqNkqQ7WPNlNWqEzr2ij81nmqCRY/4PvPr8ABQcpWgBOWT778B5
mxaCrQu3AYHTQEHPAU/5FLU84bYXJ/rzXNuWqO/dWgvYZwLrtlCyipZ4CWO+GH2DZYwRRRHYXid1
oLJA968KP35IwImXgJq9rrDMwl/BekckwhCSPnJC+XEVjRTv7pbjGoUUwJZlIJ5qz10SWUsOiDYK
3SG9yXzedMeD9IDxcvvcZTFKDb2CjARpf7W/eB6MgbU1DWv4iWmoiPQ9XVRuyiOCT3EDrAcc132Z
wUyfgbiRMd7l6DYfaQVRj/dhz8rNXAep2zmR4bzwmTRn5mwG9UT/OIGTEvUIi19fnmpdhdekCYwp
FMftMncYHc7esxtf3qTq039BMbajs6FRRHl7wR6G2NBlPAKmK14H2iQyahRVa+dk2bkUbVD222uj
wURSEPT9uHJeEeyKVvULUR2UynXSPQj3bWealEZWcaI06PiaoGphDA2LFYukEhKV3vpvk9rCjWm9
rL6m4j+6EAz9e5Zi9yuCdvnAt1xDN31nqaQMHIZj2okAvkHD1HvWCROk20TMO31o2HJL831mTYuJ
O7ATsATCb2AwB7291GlPOKOzGs4BJBVs5PiJ+aPfCu0SinE3M62PHpMiLxh2D2EQSicRDYgggvT1
wj8QE/fo5sRbhx1F+Jk5ocDDApDuehOgRJyDn8jE64wqTTImj6SzbLpAlXPb3/ZMoTa92ZYk2JCx
RvcGDtwdfdtz4v+1FvgoHxbwIwEFoP54seAmi8zizMVZ5HdS1GDDoA6zFpM8mp43Hl8zB4xkDmLX
E8FUk+Vr01/RNlmDAKkWUe+qxEk2AV2sxE4SouVyPtTwfDTboqhjkq7EI+Aakdi+WWF2KdorUSFV
DXKHUV/8d4rLzBpWEf3FOjp8sGl6a9d4e4QuzuE5rvgxab98qmdIeY23wlUypCDKsghpqBuKv4Ez
AZA1EIUTIsZP4uuMlwyiUmviU11dXAKxD94lbGy/y1DlRh6tTXmnYeh4h5M7NO37mkjyJoeh+nCZ
yn84d0lV/L5goMVLKUsA18inEfJSe54qjVqFY96g23jDn4bTNqRvne8W/DWfsH9w6eyDXqseWIHz
XLvotW5lwLEFuzmMo5vkKKnVPuPOQU/se/AZd+hFBuklke5oOyNVgzrmOkrpqsPjgR1ct8Hlet9r
/91m41jOXHfplPNf81ltTa3Tyl+RKLsrXMmWMxRqW5mMsf6aiBBufNKydH3zzO7mMUoAgnn+y9b/
ELQGvkL5l+dE3kYH2CvC0ITr1gbCSvfxU9YzVe89j8ycn5b0MRAd4Yz1pTXIVhjjes4i7D1IFhNb
WwAbQMtc6fIm2kg/RdxH/lFJNI6kVHaR1K7XQkMTD6gtDbPPJfO+Dx9DIBQaz3Awfdh2EMiE7MsA
dufS11wJM2c3pfw7vSj9nPDpb8/rJRZfkcy+oJMQ2cAcMmyBy6qcfGdVVnxuzCONkhxGTEB3x79w
rx3KWEcavPLazP5UJkU7QD6lnMSaOXXun59PHmZnmbDYrTb+LgQYUgcRQIuPx23x+reS/vZrcmHT
DNrW6KVo1G+Rb3rN9ktQSh6MssIqFiXaqClbGJVuvHKlyRA9IN+NeVzf4hRZj/i4XN/0mL5O3em/
c0WleM1Q7KM65RdZ5XazHnlphG4uGxN5DsGF1Q5lOQwwkgUgPKWITvqcaf7yJghigBZwl13pCtBs
SnBVr4B2FvvpQVbYpjryr+iDOL73+uCuMKFUock7S92gebW/2ylSdPx7JDkqRNvhFrSoFx2Wwudv
ZlRs5MOBYb/+LH5DTw7yDovWd5HBMD9uFcP/IZV+1HaW55U8xVjoy8nOGOH/3dh++dY44qfhWxJV
K2bdlnsllsbCgz/8C8froSQPN+666f8m+62GfgtXmRW8MFgLY6xxeVmw8SkLQ3mPYTaJij7Dq/S8
mntti4DQpwXy7Fhna+aotP7bOxm5xiFaW/kxaHlprqeL4vjZdkOPC19EE9GKsNT9kwBqMb0osF//
BysecR5ZzA3iLStY3p6D8Jv3N8543/SeHFwicWN2OP/n3DkZp1yhCiJNmSkwk6LcG6iCxX8OoNLM
uj/3CR/oOiiYrYSSm9WIEu0ipskNf+QKUDFPUS81mKfW3AEMA4pVFho14fnBhqzoF1xvuzN0WezT
rq6jFe7JQXXyXvF3ZdNw9UxC8fo5QNa1ezyBqDu0WR2VUnStziUhQBt0ZcORKutlpsL/zESi0ppF
QTAslxkCcloYdw0P/HQpdyRQABvukif2v1/+7EscRMQp3KfwlWbFeDvVS70HER5spCIkv+W05W3K
+veWNIv3kHaRfBRQbO1XjZjdPPQ0L78/EG7Cu6mzRyr1obegbaHPQ+vxIidU/c5/2HcEZ1HpWw6G
Cd3wgOAA3OXgIu78nHYpBYmJJW2l+Ci6as+NtLyZgdVAS90oL3ZHZxz4GxM3IpOoojoyHlR8p7V6
cQ+v469c4BQQR5xc178g7236Ln68qNYGkn6g9PMxkcj39bgfxHcoqBdBa2VfgjHarDR2kUeJqXb4
hSPVow5ruZO6PEgiwvEGrSP07WycN0GUcp3n3UJB+Bq1PFbEn4qsqv5QhwXn6upyffN3kOwY7/HX
MjGK+efZzwFH0tJBrvfuOXUYJ5z2WOxSFiTVQUwI/z0zmQpwcGf6EGY9uRBFsYunK0k8PF+Y/E3B
ZjBXjZBIOQjDU66W9A78jcqymum15w8q/CpvQe6vsnxt/yY7scyXBvJ68UVjrLNkppG/qX7Dc1uX
xfJoEpmFmFvaGIwSdqp4ymRpEdkbpEoUEITpQD3kyj0q6cHSeUfWN9bV6iCK7Lm51GGjQJRp7hmR
8oAHQSEpaGuiOjAHT1/cXD8d/YuW0v/ZD9SyjuIPPMw7SZipoFzPtO4ApZ3gOe8Y2lJIU9qgYn42
J0FJ0xMlVqeIZKRWgYqMsts5IRXN1B8L0Bttt5FZ7Yg1QoYOL0s0We8KwmPbndLBSVdb9Tg5ASZR
LwiEbDXpSdvZ/PyxFplx8FZMTlmqPDoTHYyA71CABXUEi0ZBqkCo6lS6SLztXpMLXqSmUkOq4FqN
v004pFd8qigRI+35KAtu8OPKgtumV3tcx9CVjb7cWnsnzx55eseAu5+XrJUsDBsAkK/xmmTT3vWy
NnBo7BQbv8iX3c304mwsli2eU1/IfpTU6AL5SvlW5PRWRdcZ78U3aKJoHP4rieEHuMnov+hGAk/Q
4KOykC9rybXipLBCqHqMcik3cf0RFm5SypmLrTthyHYp9+BRSG36cNvmmImipUhWZpVD5EnntVua
muoLarU7s/THhhOmm+mkzVZ5aMTPdjYXztKv6hCVAYm1HaxFb7Cmquk0+Q52KM24Fcsa+XmFpg3z
9Iz5yQodNSkLnQ/hE3DB/yi4hjLe98enTGQAKrGuD7CnMft3rULAXksuXypjVMRMczQWQejD7wyq
vozLkBYINaGeKuwQlg1Adv4X/bzjRyAuGOYSm+/iM8eVEmOLcF08Vu3b+yFYr8/islAqEO2CUUBt
ilGmhOzdCZ3NxwPjcrSK7GoQlE/jw2mJHXln9BCTT6DO0BpN3kXPUeHjIiEicJNQhGHCJDJf7vAw
CJieWbrZoOoIPcYBCXq5o0pcWYRfqSBTXKr0+LBJZzT1zy1TGCySec9VGFJDVpBD2F6qf3PZBXR9
VAFCqEURvcv9UXWzcbW0SXL+91JJv2yQeWCWAxmaOBjuwrGWi53/QJFgez8VznRCruLEmWvwMiKz
1M1nGkPo00D7F6KNFoPjp6/VdwFQMN9QEo3ZLEUPk0CcvSO8XKCVfLdXWTpFTwTJ19h7G3EY2ymG
LSYbgIapURWyk5MrWYQUPDsEkrEG0cunNQpvjlrc+vNLOGf9vXJV5/dgOdLkibyg0/e0Dfyc31+l
uloXcEQDdmWn13+02zKatucSI5lKtos79otSXwbs/W3p46g2hfs4gCNRoQThqUuIFAopt/9LpX/C
GDjBATzIW0ML2kuMuxtp5W5SPJAd805lDRJ//6TN1BcYafkUdQ3/P5gnPjf9+5e9gZkq3MYHV0bA
Z+sKglKzsSfWOCo4jrDXgu2jc82hNNePddeQkUJyH/ILGADMie1Mr3kO3DbVKlrypZY/K5A7XIkm
ZgqTsXeYvFsO/viqq+gtuR2EimPmzgPKQ+NxLamyfTx6SEBwgva8MhirP7SVtW+UbUV+GvNmHINX
fgOy3OdcfdelgnKVX2VLPQTvyz8xsUKR2Qgahs+4z5iGvF1j4nX5ns9xKmP924IeUk0fI2ypf7Io
RoIgJSok5xBg/X2XhzfcBTqdSladQkaHm5KyqZEyl26k4LePWamOPaBEaa9g+zoNV2eZcf1s8XGB
AQPBnOerZkxG/B7aGyHY1jEwTrZIQ0Hb4FwU6MfJYpzpN9nKWlEf9m7udHwJfWy7xlUeNtC38TDX
2oEJLaA6LJxTO5YiPoN3pNN/MfcRcfOk+VIdOIGTfsCajjShB5Qki10B2wMNTjpm/NiNEJX/FUxX
R05vWFWoHoEDI7+g/YVZ4Viiq9axg4eE4qlQeISDgbyXqMKWUW6Q/pZXKfHhV/omh9GH/rmk09A0
gHVDiVpuv0Yd1GTDtzNeQpLQgZ2OqgmXxrznfbU2efvtfzbO4pzuUhEYwgNaUYN4eOAN3ju7nvZd
GfCkEn4g4MCJEXpLIMLV8wY4amzbqeTCzOt6h6G9ZDG55KOc9dOjiIe/ep37LMu8zHOxuHitHhM6
i4J1KfSSO/PTiQRBXMj4WhsOfQcXccNYZCKfTFFG0WncZYDwD1rEk9jEjeEa1/gBOsUF5/2QPJG4
oKqTxZ3h3iKeseqiKXeyR/MjZE9LO+4JbDv/5Yah+cnuXg9NmIzPZSjNfXnVETivZ3JOCwGNWFyR
bUjKbk5HcL7PAfYd27Gd1JZOlh3YpgQtWxBJCKkQkuf+E4Q0ZTfu4uuGCkUOneiDV5sKrvtxkFxx
8Y8IcSavcecr0F+43z6h1IH9nhL1HzTaU+EIu7tukZxXH1Oaf17tSgdSUUQ6wNYs4W1a5/r471yh
78n/eqn0nkeymiZMX6yqlT95pLdgxK7jhcMlzf1gocVFQLVuxfVpP6NJbRAqRgqJ4DiOBwKVhrvq
OyBEHR5WC+Gc+I5Wl/kt6RlGKIbL0G+MEOtkYLBsxjF4lgDhY3zgORLanROxUvyUlJ9iXJCcL8QX
FfukT+klwLyTOgo3e8H4WDYct6wDGEMksThaYHzhi6juL4cM9TEA+zoYkx45R804O6dd3ZyII7P8
riREMncNkCzaMcJg0u705spehbYNvur8I1unczbgLXbTB6ob9mkgdfUapnz26g/ugICrMwFwVGtX
cPNItHz/2RoRltu8jK7AhtdOkaCnQvUMS3vUaOVbRU+YmM4Y03ymLtCaYwqIatEquNgpr5oo4LC8
BFfAROQq+QKIlOYzf7UFP2YoOf5zFdVhV0h2lfbscACA1jt8J+Mev0A7IHXdUHEvuKahHeZjq7uO
3+q6gC/cqLRfTiUKMb/WuFTMTOcLkMg9M4yFoOQjbwj6t1C7O5yXNXXDRb3sDBPyDMMDWhm9G8px
0nZh6+yH4mBHRQImY2H4gL2gizm/cWngPJdLp2cgvL+fdhQ0YTeEpRya8MxWoS8wa1eVvkoOJ6BV
YTBkjm3gYjhDyybFqCrqFb0S/AW+ZC6ClYrjvTVxApcIZtwMQIQHWoKLXYT9u5aFvL49vdCoZ5X3
hk6wrfHcp3KzGh8Ep1YJcNI87w7ZgPbFS4qGyM0WA27BWUbcVDgCkEw0Zb6WIfX0Tzd3isGfk8mJ
sbJxpJoiDY/8yTXCIFdokutEdTmnGodkl4QEV0yL1elp5+pVNxE+XGGILMbEGKL+kwqKaI1X0igF
gfp2UTsIWMGLP7ZsVMWheQBPynAHpxXWIS+gCcoB/9+aOiaEnIlXxAYMYxmGSlD6TKimSnsMYHSX
6mxsMztBc1T6q3G/Dgu1ML+dof+dazfHb/bX7cC79mGBBPLaaCdfGLCojVBwYTMORUzGbg/Q0RLk
znz/c8G2yXmC50qLsGgHbdVrqfZw5keI9Cgjr/ErG2ZEHG8cfpuqs2z5zi4hM4L9JQGpz/Vg8C24
lY+5LTeR31BdZBun+8cB+o1TZ+OjFmNHtWvzBt/8V5bGaML+32mYLRa/vrM+63+ptxpBLdPZWng4
eSjRJGO5JEWy3j9ymT1S2t2LWNGd+RElUBlrrBDDQq10cMn33eyK9YclHil1QNNgItBHtKMfPdUc
Z18pG/TYfP7XDpN7cOW5rwkSkZL4FKYwMIQWr/Ym5CoV2s/5e8CKv/fYuf6U9YiJe9KhriqqBDQR
s38x2ga/9kLNm447I4Vl+rgwY/ddSLvejscgjV2ZqiGPthnTPmvBI80GSzRz3ygsATi+nuWhfxOD
/irDKJFlLnzWYbQeT3m1PUZWMe/tO1ZNs4A9Teb7+Ohykz2QJZOLX70nLuwVj8mKZYQrdianpi1E
iGWNZdOZ4Lov8ifCdhHLAnSel0XlRayvPpsDrUbMKvfsteIkl1RAid86yi2ht4I1BQeOqjA8RODK
QiGGzxm1sfEgedIGpspPHZo6n1yBBbTfkru5/6oTPJG7z68OBurhDDPU07u2thsFFp8jjnZJtAFF
5nQU9q+oaPsCrmbfs2twhdvt1AdQoxH+IK6RNoQCVwSTl8IX2nZ1o2gtzPpV/srB05Io5l+z3oUD
pwGJUl+KoI8Dz6z6xgVNvYIJeUT348UR9WxxOtdqjod0pXLUUqI/Yg1+EIbcKbMcxN1Dv+0Lm44I
kkVuceONMoUo+SdfUCHwPgM4kfM6mZfSSZN2TthRa+Ut8+eC6RUrsOEgiOo6tK8BKdhetJYE2Ojd
WMpFY0gRPryRj0MP50sYVfC1ldv38vr7VFSSA5i/vY4oV4pXf3mhNH7m1pB71fVLzfvtqSGvS8/w
Cliunj3UcglxanML35t/yQxp4ll6YJxCCnBkwi9BovFAwxNVQgwZMdGdRRxLTVy6COOLRwrcfudl
CMsLxXMjrddSLvCsfYgdKXRo0J0Jby4dvFN0OrZVL5wQpEXmSvV+banfZKAovF4ttFtjYZm732W3
lstq3qhXCq4VBaM/vORXZVUzhbwqIYiT3rKxPS1rYV0IRJFQL4j3eJYDkTfbdV6ZLDJql3SSJ1D5
vd9TTqHEdrqW8w7OC1QG+hsW1wqz1egk0UHeF41jWYyqLDDeemjaV46/qheuN1lyyyXr8v6WJWZX
ASqN5J1on3tYLp8iyUVx+a79jvLAVkbHop6m3dZi3lQNIBjYLfwIv9L7WfY5VUzMu1YfsmoRiV52
RVAyC0R9GKowkpbizKi8hvgfmEqcWDjsdQs3lSaZbuZqcdVHJJpJdbHZPok8i3yid4vjEafbMrh+
mk7TCCtq+Y2uWYNo+tyv1pZ/Djwrz+3q4/vOY3FI/QP9Xfi6SZp+gF9SJMMeCYPtf/qOHAqyr5Wi
2pHgW+ASBelDfuNRgRBCQ7pkD1JLIVcs7rSyL5SzaBQJtVd/YHtYB93QBoWfhR+tauHzDuUUQqCr
IJBd+JbCEcz5DmiBS6vAdHi5GKZFc/yLMcrp5wq6Dy84qO39V/duXSriXtUgdg3aVsRRVJUbikT6
2dMMCf794oYwdIakEPtk7i01DpHY36OnNY7l0tj8cdv9cD6Q9NRl/Ima47lbleSaDvk1+xyndnuj
53LWPmAoFydWDueiZ8yYbHL7E6fQkFItGnSCUQTzhI6X4Ip47sQXCri1FO12lP7WeIBrekQ5HHEF
LxaUJuioPGYer0bfxYdDvTO+yukdDhKR1L2hc9PnFcdJ70ZAytu623XUdDODplGy7n2kvTMcY18A
wdnwYcW6ioJmsV4xI/ZMIqgcNUK3s2ofH4sbQOqlPDJpl2U8IeFNe78Edlr7st7R2UHHCs40Poom
HkxKzbvkywrGADN2m16NEqCK3lOP9BXBTFlpHTaIClR9YzoYSpbIV7mloFM0od2MhtkeXik9rKSo
gedy57iFyDZfKZPMCfVEM3eZxjiBUOopAjGbo4LXs3O8czGaC7mukI9jwjiRt/SUuqoTmT5Jw/TZ
WaS7KydFJLR/Pk1nhnWyDuUE0u0tRiQPdLyVlwJCst7FbTb6z9KLrXWmLbytyHunFRsjgn1Wy/Bj
ZYKhqmSc+OmU2ZriwMQ+Y9crLuchXwKKR3jzbJZZX136Sr2ux7RMA9KTlf7Rlcd5cz7nGFpePcfy
SPpEYapovvefsECTiROQcJyX5R4GNmQhqvgzWbVvks35gZf1iJc9CaTeBuIbWqWnr0KiHY1spqtV
H6IWzOqHzSB8mVUKvSF/u846GZ+2GJ0ZBTfBJyc50ePM9hhgDNG6KDUNUpUGumk/aZt5KjKrbXZ2
TQnalZ40f6edgA2V6RTqlVdrbd99xyPjT2OjxbizDpUtGuOkF/fGjHQm2E1WXVwbB8o01HF5uikO
GqiOxtsFFD1nQ+WZU0RIGb6z7c/YIEr0fKuVRBJLLyvohITsymRcyaWH0FAvGfG48WTvO7RDKRmX
krDqF+XuqwXfpTM71xoESZmGFKtjN90xwJihoDM/3qhB5sSN2KBJOtCE+OG8uLCr4f/UGlohjO4l
KVWmfl8Uwugz2QlVG9v5ObUVmfyzE/h9PWp3fmrrrzoLI3JRnijr0SfyhtiCyj2NT+or42mase8H
FX6d0lEYE/kuy+3Q7AV1FdFbfj3cEG54jiHgl86J70T4Xz9+95E75GOzPXE14ma4HONOgU7tZ+T/
orgiQ/R4XaQkGYCvebI5BubTJIlwy9fYHejPwx76joNAPYWDqhosIfYIGqL+cGU0wECxm+abnH2Q
rPPrPvuP71PG/q5wovPq3Grwxe8i48D1wC0rp/j39YMumo2lCuafVys9bgFm1sfeg+DTMhxiFbCN
rHhrWyDXvIxe+1Qgjjt3s4K6SYqzwAo/KsVeIPJxo38ml8N7y8GsbC9JzrZtk4EmAuj/jD3pzE/n
5Oqjii+88uM2FB/coJeiLiQXOvv/bdYiJJmv/frZNWR0k9/TNLsAPZ25cqtaW3m2NZsj9DPM0GkR
zpo3LpCkYeNpejT/Dv1tkZK9LMIxJvjNP+z+Pcjf6nV10SEeruvnMGtybiZHQ7UJCiWA82hxrXt+
SHYOo1FN4Xu4RNAN0dfvPlkXETvcK5/XPDIHiTkxwwOdYFOraDwfXc7aNmSQ3Fp1oDokEeNqVSLN
pz1JKagsUMFnXfKo3xU8owFk31+XIw7Q7QqErZ9VtJQyTC1BYm4VIxf3CfMLiqoz4NjHlZfEtdt9
uV1o0D1j+7tcFAK1iXv81UupFAoEZfGVQR4QmP1y/RizW4PmaJBJQQdHKpDYsTTiGoL9jRCoDifb
CP3aFN5+qFL0LpQyocLDgy5JJ7PUpyvNVKRE2lI/lpQdr2nCO0VzqzVIp5Ur0e5MlKwJYdGnsdzs
iP4ToBh658k+1+1xYsvrg5vrezouSvNVeq3PDPSfGwFzimr5BWluqk1iGakpodepp+y7vcrMabxT
OtP7a6LJBtF88AWvn+vhgzdo6BeTBwK0ODN0x7WwG/goUTLH9eT7OlHlvSHuZ20GenvVdn7FZrNe
+nn7l0r5m5YBZsE4z28xGFWdfQ+8KCUToLYSyV76qSsPSMmSDm3PIYpjScuEtbtfBQzHIw/Ob3CK
lu1WXi1B9TKDrflHNlykW7bScazVTZ7+VkW4nL62haHQHUqO5qmT30sJYCYmYV4HxrKHnUKcJIXw
OEky1qiqvRNyOcKRNjQQOTJee04+6RThuiz3chRW6PKJZGXsu1msT+HvSIBjIX+FDIcATs8/DXJp
vzzjgg0Na8Cs9i6FXsP8AnUez3lFbYEqJtd/t4FNkTMkAzld/ryHtjwoknSiygzi7C1FWhS3fYov
S9IUe92oaAd92F/piWliELPa+DAlCFUNGf+13Ev6w0+iU7rYyU+uApeysz6Ug4vCl0oNAwG6pe98
FhgtVjnAU6l5+rTpoV3ee/BPpWu/Sx7/Fn9PMstBmAyu1qiw+PpTclJFxAo/nMOQIJA0Qa7GEM9Q
WJo0Uv2y4oG4RFGoZ0AMXoRw9x4u50akvGsLgiNA6DjMWn+UPYt6UbRMx74FPlGLlZScVqLxXMXe
OdsDirc0zJq7zyoMc8yEBgdDOr4pI+vepj8+T0OufqhlNgzxMW6g7o8IjYj0Nc/IUfY6zM2n3qZ1
T3b60CqZwgU9flxCpiXV1ne4TyORVcp1M0oTAk2BBZi9U/xBi9NkH+B7fZiqWGCXU1PCLws9GZTE
IvgQdX3W/+9GD1Y+qZXpe7uMx6brOIKFo3k2fIjvhVnrnY/PNY+Jq99Q7utqAJIcth0vFAeWpQqv
LuuqFEGaOyAneNhOfWZdU7WFy8lQvpRUyba54UqWl4cM0V1aR+fuVC2j3HohYhCu6pou6tprhkDb
L11sr5quKmpwgLG8OoIh6zJbA3wX+OGyUo+ppPkTXV/6g8k8PTr+/xJnACXDsUu1qQr8GL5cSGKJ
9DJso3NkojVT1QbHJDZUNgwPZgU0Tp4xDVe3UHFVcObYoReSMTtiXrO0XZkPmCqqlsMeAK1o0UDo
G4H1FLmAGp6B+NS5MfM02VjMn2NuqFY1fpAyz3Bf1vfBMpfKaDPmjSVxt8LTycvhqM8pWyg9m66R
XEb0LgS+gRneBFMYNf8YP0vnJEZtFrwRbVDBIIWDqzi4xSUa3WPfSyNxg0yW8+D697zMuiMXfN4I
k7cisvhy4tenuRiDSKJPM/5/oLYIcS5toMLYZHYQohP1QPZxoDIGlM0FSdFTosM9ZDM2a3uTe7rw
NvydCFEHFskO4FKlk1XRqXZqZn9JZ2hdvXmBgsWwWIkjnR4PU1CDcDevEod/1/3lvxKKUEvQEoBx
V/c95Rc8y+8KPXPN7C6YZ/U6Fnj/LmFbmo+zz1l2hyY6g6nSMdN/p5or3Uao8xKul5SISditBzHU
0wUwyu8r3GP9YkgmXk8mgny8vkX4YlyvbOl3e/of+Lw3Rj5GPk2O0MTu6phD6uSt5RXmI+GsGnS2
77XKoiYb4NOwq6c4KW9HZMGu1khzJFPZirF2k9GKi4dGWWPGkxbLRGmv4KiD+43QaYRHcSlWyISk
7YqR/LxXu62s9b92lNEYdsBK80fpahkcA4hdGKDZem7Ce80jTVbmcMseOMIa/UM5UvMIWngc0qVO
1C1alOEN55/66BPnoaI2icVqrr9YyR6zWKzjOPuVLFN7EHiw7BUR2TP9tibvNCxJsEWKVyuAe73V
Nfuau+SBQRB/oc9odjcLs5sihU/ZNjR2TgxG0nbKfYjbkSkHVpaY35IVw28oIROcNB7OE3slQRYb
CtGdV4bGvnBJ05MB+eJPMPvWFzQ+gZLRYCnIsEo7RZzWrKvMj4Q1w8rRHUx+O0qfQ0NxuFm2zY3m
+KOkrNaclAjho31xhNno3GO7tuFcIw8baYMUpUqw/JdGZOeBwY2mkG4Abo/Y+hqXB7ASBrVYXI5o
oR99nBQe1BRygSY79OKzm8R38GbrYiTwda7XXnnsz0wRK55Mf3wN565QWWV7v3+eG5l+7bmgPO96
2RwIlQdAPZ5Wc+tfUHg6A2Mc9LPmhMj13FegVZyi9r7MXg9or6U1X/2h3jt/HSdzPrxXQHWTc/Ej
GujdJP/RK7JVrT0hfh5zEVWvaZ6wHXcukXxZyZHuiEFh1m5ugHyZXT+vaBS1aV1JC9BjEd4Oiqta
upSHAjXaAuPeUe1fWFmsvOReZiWOAzmZyIHNp/rARIhNxdrgUQwdxKsUtUxc+YAnHiVH/1Fs5+OA
FZO1x1dnDHwgEA5MSidrexOqzhAVe+3g2FWH1zM4+zh0QmGbLmaQTsSbAw84pSR044Qp838M8nXz
TtB7Oj0j9+Ab9ETvPai4ikQ+2XlwYp85LU6db7jBFwzuIHc7XsCqVAAH4yFYgWIH0fnDMxV+RqxG
AzOIWW1pSkb3JFJxQzDfuWkxD6jOyQ1AbdxuhM08gbuDSVSGoiK4h7BZnjRyoCjjTirjP04DmG+t
X/Ls3hUArQBB/pFXqUbnJHQcvXUqiEx6SubYafUxfKN74Xpf661UvNUSn2sn1T4cWlaE8oPVTVYn
+LioncZvzf/LyuU9NKW+jagDGbO7u9PQTn/+3hr8aSalVm2/mlg/eXZ7WpazKrwYbfplqThQUlto
Hxl6Y3VdhGdxIZgHl0gpPiSfbbr4MAV9FN5atkE2DRHVmC/VKTqVy7FXhJ4Q77v9H8VFbMCCHRH2
8OWJ6pGaiPvO8kHU9fsqcUIKY+bLJreBskHDBKvdxZAI6f2qcGjjkBEHhJJDBAF7OTvkUoVhFK5j
y+n7fDv50pYFYR8qWsQvLDs0ojOxgWVhOBNd5xsAlXUcoWq6JTqNF7RbMzA7iMO7jhA8+T/B//lL
7uyo7d7Q4qfCkSUfwpX3ZyCL/m9imrAZfFE/hCLXQ94N03FnKWOKa9ZrpAP552I2XA/nZ2dgb7Si
IkqaBq4pD3Kietdd1ccbpuOPM9+rUtrdTxYqHivTQDqyv68g9dR8F8ZhmnturvHvmw1tg6rOLyFP
m0ZxKSFqbMUmbLOuzKoh6wWLZebhJ+0C2ENMsoP0P/8rH/XjD23fW3sYnWkdDdwOuX7LX/1DN+YL
Y29DiBucB4Gtca+VSfUUQNQjlcgMPAI6lE2r028D/p3o1s+A/2GFqu55cM3CquOpdiNxFm5/jImo
iyReMjQSysbFWx7qAh2/8l0/oIYZAZi7QgqnUyHTIXa+AYmGW4aFLA2a0jeZfxVnQRedOXrlaZcV
LC0W3Mq1HUVAt/G04LvR1NTSW/JN/YKTPdOFmIEU1RePU3eJch6us3HiP4/03RxlpWvQT3AkIy5U
3xxvtRHPZizh93uONcPVThw5TPf+PiizG0oACp9UQQ/YxMEAAEoCbNxfCIZZjbBRnoNW8CiElLtJ
EHjJyG7ojJAAseSPpMehxG59bMhGgjeMg0zbvrTokLXQxejuYFAXcPhXXpGw8u7e2o4Vfk93+h/v
sZkbBonnKbVxhIpsOaefoC/y8km54VXzWnfpI0zTcxrDc0jI/qKsSYM8QE6J6s6JwWzRbFmyQoXI
XkicD0NypflkeswLTPHApCNBKBIlq/AiLLG1l5SbuUBPGBI+mzI1mqeODsFLXTZJ7O37ok3VzkZs
EPQv2YYAOCUNtxiHWxZgWQxJpElwezcb/ub49MdzdNmrgBkR5MPDfyQcz4SF6Kekp+GBTGBGbB45
rNik2M80w2kHlZNEBKpsIXGyx7qkJcIs1ihI1cclFi+hh9paWdLRhvELcqKb4i/6NkovoCJMlc8V
B1VlQdXZPuMAnhr+0bBJjKHUl9iJhvhqGF/6q2EyBo9N4Dcxn0VYyki0QuZMLi+f9Qypj1qFmnA8
ODrQHbwg9ln4H9zGLhnk/kIMzEHeBE0DgMfRJQdMU15cllLKi/Z8iOEIByV5rXhNfu0o0pO8EIYT
M9XiElPKMvCm1Xgmh7+yjky4qXpc4Iayo6uWi7booHWSmAkrqLMOYG5oLSPP0J3ksMGy4aS9fo/F
/zH7jRtMIZw2B9VGMjxaDN0x010sLvqPsIs1dxhneantfPmvpSwLBCVTu9/dgub39RejKqgOjcGY
DyuiCEZPNZTGTXB4EEfVFgt5/AKvFvL54WQOXc4leziJWnbTs7FWZKOeIka7qnnxfy2+rlw6Se5o
vKEiVo1iKH8NYvK9lPvsTxIlvXHLQXB5xRzctC6HLWDoNCEW24ixK0XD+Y8CZK1Gr1KY7DL/+uEp
pgcGMgnpfmO3aCqP5/47Li781VOQdBYuYacew6OE1p/jpWIUS4giT3VcEPsmpZQ+9h6F2xeEbLIB
XD55kiOOe2JwjZYQYDg2ps1O0Z3ZaaZqbosvWJkZUk5CVAjwxY+xziXVfpiFWjh7JPo7KDciWsiM
GMaaWZclD2pXrz10KgWhjxOg/Ua6HDZtAfOUi29/Gq0JPxPrOfIcs+qO1axxIVHFzFmX+AsHVGRv
BqSceAai99gX+VT0akcCHfkdLZcwnBe0oaha1EImZbHErM/ydilgvApbieHAhUtTnjSkrbWTZX3Q
piXLOKw00I8W45twQS39sC/C6Ms3FmenaP+nd3zGP+0I1Qt3HEI+COviYmE6bR35rw8XvBTjVwcK
trXDGlBTq8drzN6lK6gLnNOi0j2OQnYtrGmt6gWDMw+izkokT/eGf4KmhXBJYehF56PYfTJ0VQZm
JJjlcYEhtFmxrhm1M90TTcs9Zn6+o5OmaTvIJin25kRSv/R7yzrK8q/27RG503ITqawkxOb4jYIw
DgpphpLHllZPVaWvZATgCjCnaDhE1gc8aI7HUlzppQs4pggak6/imh5ZjnIYRR1U6fIGSleLbPHq
gNa62rt/Usoa9nPq/jHCd4EwO+V8VOUd/BDOHfbU6YVqCt+G9T5AveMeSNwfgaZhftTCbU/vilPG
ySgVgu0KxBVS/Oxzkl4ndeQnyJiFHxt9qvMA53ZDJDZkH/EYEDcRgs9OG3DKWWAGTXa2TZTbFhXY
QJR1lI+uraZxuYMb8cRWMQlpsidzaBtQBi7YENtgVfze48Cpc6ksQgnQOIn7vGoV+Z889iBXog0Z
ITjF8MOOi5u9KCnf01AXqboiBAk8AtAGkPM2IuUGyorFz87s1v8UNMVT0rgBmlooSwb4wi0gA80p
6AYnTfYuUEysY3CocFwmQS6DcNNFZiOZ6gl5xHgESf2n8BsLvObYHvLVYiHVoFiQZwxJvSUHmqwb
hX5qdocRes7YDr7Syz9WULt0KsSqNdf7n5f+I29rWvADCn9FniGkZbeMoNlEK6mVFzD7WXrBCpdQ
2dxwWqRAa2wVcJIqUSWRSSNi0AmflxCQI9c/njxWCNW3wgXtPwLaheYZQ3sKyH/AxLJ1GX6qIb1f
1kJs7HV3cqo9m/w3GsTIuBw21c82VQPDlqPtllAKCm6d4XhF3gx/Jr+5SowoPqf3T7Oi7oOYWPm8
a3Ctqp2IruxuY81Y6YDP0pd6YLhGCg8qpkZrO8LmEAxGZmVPdVu641+L+DsJPklCaWP0afoF7GnX
Qol0jv+TcOJ1oD2+Cr8XHXg0H42JGb0TnS7LOw09pLPN9qYwaUDsOZwqB4WQ+j+ZptfWN4eaqj9y
AmaobRHp7kMAEwNBXB2T4pouH41XJ1Tv6EepbZOqX/IoIFkwgm2mDaY2Zbkw5bHo0f51NKMgIwmm
fxJyj5GcLnmFEJwQDRd8jA6zalISTjdVgZ6BqpvthyO+A+CFkGxSPC5PIEzl7HsOTFMEcodUycL9
zVxEJYf5fxNZl/vLbk+3MnS5Na3GHCv4fo1/xYI/FBTndJKstpLW3y4k5vUlq0VNlI7tVEL1O81n
sB9h+9Q2t0U7+XSP2coR+tftFGw7qkjUyMfQj/+HjYJrh+ufovWVInDKiT+xYpbhQR161v6LSFpy
mJiSFAmuyobEjjMADi3yCLTpRh/77SBHK7igy0p/XzJDDbP30RBhUq75caE79NUQk0AiaH7HWJyC
G1zdeC3PI3xy4rcoTwZJT9bKJWAmxyG1dHhNzEYDyrJYJBWDyW6W6a4WXYCDrDgrDvgyKFk1DT4l
8oPIgrTlDSava5/iJcwA369UipBndC1Qzk08dQYsqiGNSlvE8ZiZPNrndBDhR2RdcsRhmNwmPMv6
RlvkVH/YCaZVMOS6sn4B6YrjR2HvFM5HjPbdKl4BbkReTq9dpW+c9m8UoIImOu6uNB87a9xW67U3
951EQds3o3EB+AGyKwNgUHLrQKL/+8zqdhxPa4U3RjPhTtjZQNLrZPOqF0mRx6G7RkHTWczCtCvE
VB1t1yajc2dQZM5jMbvMzDcmRFFBAhhWh2mjmISLWQz/W0vSbOAnbmMH6Jwi0J7m9tm0yw/GZhm6
2diR60JtOvup5bkuSeayFdmXLMFdE0o6wC6FjMeO5qfq+hukij2N68iNnGkuDcpLm6RqONLR9KW7
A0vqztqqJGb8BuT9J5Bx/qjkd5Fdpe8Iwa+MQd4pmnNWrjjp9ZOu3nNNp8bKzIGIdJeOzvYcXnzo
Icpx2JipXFsPrvqCWDCW2tTAE398SBYgl5+ZcxpL/1Agen+6XFbVJsKyrQV1oZH6DepVg7ySQyGf
rvJsQ1sXQhd35yScA8Gx2gtmqmg1qxTFVIiYw6lw7iQ+Lto4KZO+3pPE/rJB2+ZWWHvuAqhl+gpg
Hu0HVgy5xNt4U3CHB/+KoU33Bi6tZh89Y4eDvWXkxsUiiLA0BZxItlcvfEz497Knwc1c66gyCcjV
Ewoo8dJo8n/ixB7wvuStglWvyzTVRWw7QZuBivPaB0s1/c8LxLeFlk4DTbiR0+yp+kCU4lmQS+Ou
kYaytJfJvAvhA9+WBlMKjbHvorxm3d+ib2j67UhGgIGy6Clz9q+U5q51iJNwvUU6oZqbFzS9Ov1K
sqJY3RTyM2nYKUMbZUOJIaQGvrLHTTPf+jTBIaJb3dESyp+xu4rVEpVjboxsjI5u2/8cioGRTfwP
RkHIH9sw6upVbHWrlAAo7CpIxlG0FdwoRMfQA83Pjb+odPVScyKC0ETrFa6vUU0al/ywwKaojbIk
+y07GaUzu7xeCkRvdh9DB/UdTP2xoLZ7/DXjUIKFa5mbeVYDA106h0XvOv43z7AA7EPvDKrjeuxC
RYQu4Y2QFHpllGwQOtiYEIqo8rpnharwIBZkr1PPrCQNgK8b05qiXGGLcIw4C9iaCFOr8nfU1sP9
atpLsGQTZdKH9CyuIBBuBFasOdsffD4ZAHnNZXLxOily7w/YoDykKwSSg8Nz1NC9htSShJ15+Taf
lDbFeGQ3gvLZMVUBgFLY/2F5zKwYGEQ0ieVvUCn0Q44xN6EBWc3cFu4G1v+yQY9yQamxom7cqVa8
FDYDvO5vlgD5EES6z61e2sZJ56OquDI1Vv1UPZ3/wARphfcnKVKen1fpCEN1PTMgRqjCzckuA/FK
pMVo7Rf0cWbNzuv5M4u66bR/Q5OOZfXQLwhGR91N26ku45J956XDNDJq14iQkjWTFJxjiId3kIi7
N9WMVny0CLikqyfHDg9XBA68h2sXFcxPMZuyu9jN86LhH9jOpkNAaAk5Y26wg38cVvJW92vPVAXz
zuK497Xm3ERcDDhfDKs2gGnduzmAdcGI+zqJLLjOQqpGlY03NJND+vmgTOclcnWDYrf30TNeajA5
wiGgoB2t1cdUL6mlY2rirjCMsjeZUhTu/qD4Jpl7WOTmQd+Uv5ZJX8UPCaCwERlq5YzR9DlqanPc
f9F7rK/zzY3ITrMwTy35VqmokvsYHrXBmN/zFkBK69WXELZyoPCrhr+SvP3X3sgcugu4DGBUdtSB
uWRv87CBwdXimEilhOtwMRND/kp7wQCFXyqPBTS0/vHM59KcxqfLlRLDmjlWjXgl7M0RCNG5wz+l
nICAMYzCttAbe0wLKayLfcVLu0m5sGERT0wn1o5D96o80krMFwzvqw8Bgetpr9qN3DNQzojMw0D9
gVS/6QW/Yt4YzLFrx+0rzU+QrXbE8WQYeM+VF5MaVk2vMDMGrteJJy6i4ZLUF2sDqiitf3Ze85LR
FPhSW9nhTQtgylaNAOIR/9wUx2Bcz1pjAi9QJWnB4cWV21sCUwCJHrhBlSunSMRcXGOzDkkVg9bU
ymXVmdlfKOoVS8tDwNU+tv6u9ZAxd4Q1JYLkE4irSXO+RAsUUimr2hgsSMeP51nu+Pn6j8C8y92k
wJklcQ2UrdRB0gr0pZJk9tfnWEDU1j7rvZCdRvDfcWJ7sJppyZYBam6b/7DwmEHjNGwitQdymvEc
s3Y3JqVVk5ZhTQpYjvSjyAzQIUNnzIrfCuAwOA/Ig2yuMskXNHHDcpEWhZwYniuC41OB+m0kGBBh
6VHbVmi3fYaGqvFXQIA4QGJ/wP4rxyjU8LtCxnNb1bvgWYKUaE7fKUlaMxt3iv0U1SsN80XESyzl
fcjq5CHY7ID3mvKXTwFLLRlIVzZLpsINvcSnBTtZRLwBGc8SebdAMNKwSWU9IinP15VqwYPXzjqi
1qrd3uHsXWHYQx1ouH10EPjJrCsu8iLfpeT1ucQlNCgcQy1RLIN8hgrMQf1QJZtp06RzBxGBTDyr
J7L+qE7VTLvjbfjeb0PvguX0pjeoJW2UmZOUSw3pQtNajJcLNhlXyJpSG7ovMTvtM1M0lTu1dqJh
wzre5dYDr9UQVzn5UGe93lrhSA0Q+8lZvSZ6oJhsloioNF6VJ69Yu7IhNtvyoxCQk8uWwrjAjbua
N9rcUdgu6HOgjLJaG1UrqK8w61+FCSodKGEhS7lOnQ6WbTs9SMuqDQlAN5ovH2e6Oko8O+Hy4keq
LIG1Yi1Qr6It6+q+IYhQ5KXGXT57s/3KVKX2uWAKiNIN8qQ5gkECNlKaAkVxXukthISdN4yGYSAb
wC2Ie61dyxTnrL2LnWo7EwvBtlcseqWkitA0i2xSsrtCuQP5s0DYz4P1W5Mr72U1BP0QMJGLBG4M
QTANBM6cUsKLDHrLq/65q2Xk1GeoZQ1X2Ux5eqZs8BrjNXnilp5a9pYnjVtNBV2sGkLj/sqYIJSe
oTmuTwHgvplOsY70q/U7lNiMe5Qhr9L6Zoc3IPyryqaLztd1NgyfdD9tREm2B/XBMlDmNi80Ia9Y
y18tTlhrvoH0zodUxHJyanGIFn+8TBST96OHuFLRX6+HBRE4jGG2EKQX+V6EfUagx4Ls9Nuxl5nN
Qy1dNRXh7YEXkOtXoo/16dyAa69ZG7IFCeuTfeyGcxslJd7g0hi9WQ+7HmXLW6AovN0u3gYn1HF5
lPpYqyKFFSwB6YyFWrNR+v/MIWejvW303wWEnR1D/lMCnIgK8FPuabZBH7Fy9RtlCnrzFpxNoRqw
Zz9jyDnTGr9yO+yjVe6OvjUqWKHsqnYHpCRwpJGvgwU/6wpYqhjHduwVHGUb889aqAxxFFY6SjMS
/Kn+dTX4Eb+qOZ1iSI+r1PEL7ldmoBUpe8DJe/HwyxGeJJn5Frcq/mAoY33tS2/Wto97RyizWUdm
zpUJJnCUDyouvqt5IjWMgR62cPZ7/F7MWXYDJkm6bMr/fh6dfh4pAXaKLye9J6fTudFlIBzVG6dd
RPjki2TtmqghlAtDXNckqWKr90jhc/zU+8Cupq8B8vHpn6C370XaUT/HTpRryXFnabH6B/dOD6OZ
AM1v/TauaEqZhqOZJoUwFUH1ty6IclW1PrTw15NqV81FymPJfLsN7lu0Cy2FdoveTblNperTFxBB
wDt4w+KX1imp68drUK8N62PEtYXzzs4ZUpQrCunlz5UyrsGTeud3PNfPxz58hVKAoJu/MrlhtpgM
jJU80wGII9VvodpKucUDgwzbKOhYQWGroid/mBnUX4yGnh1y3vTBfXl7TTgChMmsMzZ0rx2GnnfR
rCdSSeKS92yw5eBP8QbyBakcDAcNosSRKv3vRK9l+F0sA24AYHnaZESDbclR7N/Ry4Vut7k/JTCb
CW59rv53pYpQ01M1SGabrgLLM6BVqNr5BCnD7aI/eXH2gRg3V8f4gm2Ob61HBAWcqF2ySuqY4f4T
oSJvQLYiWETDzDeNx4MLokNB76EwYC2WsTjq8uxrIcOk5ftKJKyoS6O7UTogEshjeG5ZqqGAyT9E
x+0eByd7f2m6ULjaoei4tt0vYon6N+7MTO7wP0AtiLjkkM6rA0f2Hxd29IGqlgd8ukPbxSppor6u
AlK01BRVOIhT2W0PYso0MIIbdCIaWsGrhLWYvHyUWQZYT1h8GpVEukqMlfbdzthNcAz2O2dmYjXb
/ULwMBcIvNP1OK+/y9pHHf9swhzlWtc19hsIilsjELHqxkvc/EzWUpY2EBWeK05dKXS9GagJy1ml
+HEKY+h3dsAjYk/T/wztbrqF1sQP0mmtmHWlHcGjhydroGl/6siTEgwNSiYVjWN0/3iOVttHnJdn
GrQn2kBPvXS+6NODZPaa9E6P6ghqZXFEcoGpEqx9Dumfx2C9/B2cV/X9I2zz+QvioCRVnw8tA+2h
Qr1R7ZadcvKPXpnk24vFBQ5ZkP1rkQbxdoJJAmLWb/gJMNs4GRZAK1I6Dr1GEDRzcTbTCpboZJs6
4JjTAbTRIqAiMymJTGEaDHzSOYb7B9XyCMSie+U7+irIZW+tlKTU5ZzcmxI9hM3dsER2JLtQmadD
0jk53DGxfHsF8D5d1qh8byqm0k28Yp//xziWM6uqXcG9mIkCNSQ5LpNCRNPtyguPnTylj5xFA7b1
gXvRF548y5gWFN2PUtfhBJtmxk4goKTVe83Ct70ppbaBazLEcLLXT86iRqwVSQJxv3AwT4ie9jrX
HTK9ZSz4PZmlwCKziYWE7gaQyknbOqsCMsIcSAxFoI2Rt0OfBYKH4ra1zI/38HDOJ1pfaVupKOoL
89FRM5QyAGn//h91BPfRfXwcDCSHdvzT8tQvgF+Hh/W5S+lWoqg6oHPkAwZi8DOJNPqUXpHwMBjt
S7PgL2gDJ1SBsV1qvI5kzsqi43V4bTyVF+tVgKrkNDxgjHIDKzNlfs3MtZi9kfRkKIbmGUfD4fJq
6v3UgMhqNKkZe/ZRW6yGEqJI/Vz+8FVUiOxJ1LBfBy1godBjWZgzYPJXC/zhMRfaHIlWYKpAC6pe
9BE86WKbm0WPX3ZRsn9EwxqJZur7wxa218eik10SJmU2cxVvm2EotuwgMeGs51aWgGTILwECGaok
QfyB7/orCMb1PjJ5uart4sMgroZT5lYUzqORiodMQDnO0j33lTy4U3WB4LyXC9HxkwYo3LjQAigX
Npf+VmfmclXtn+yjCC1QDKrakuDoXNH7pSZaJ0A3tNass8MwBxm+b77CWFawMcEF1+Ctu9f/3kiP
3zwbSkTdjtK43lv+NooBBxIjUg0NsrZXMCzTIvfMkB9sv6Mie79mfqACaMai/DPKxy3Glx2+6BYr
mkNVMIbZBZd/rkqvhrc1ea0/GtLJKZDstGp5kxgi9k71lC+DleGsTuVz19z0doNwt+5ledikmkcQ
Y4YIIiBDqfry9OKU4kBYEm8qLjd26wdiAV6yj2zTrn70bzHaDxSwRWQ0wb+iSvnw7dmmlPsjhX1g
9KCdYdCSITcGlHqSiz2Y79loRRV29tFubkEvGWsyWyRjaH7CyOA5aD26Eew3YPZuCnsinuzNjqgx
tO73qDXz99+zSweU9QLt1enuRK7ykDzajMJm5AlfZRAzqDQSJvRuE7+iF0HylYW2FREiw6rXgP2f
yf3iBaN+sb/qafWm/dlgbWg3HbggPQfN2/FEE3hQAzwCBuBv9ArAN2pRPvuauOiiY87xjboP0MDk
VLkdlZfFiKC3ut6xxWwGWAIRpNCcecDBE+A8OH3vUXE0AU7vJgDe0iXiZbn/gdxA7dYdu62Sn6pn
jY8pCZQ8GIxK8r0y7NQHQ7uSBPBLftzHVM+g/DOAWQKbBKom+gblZunu7zKz9qMY+RDTB8bV37f3
nd1fvYJp/E04MAnFfaWQi0DOBF6OFyyCfxryt1qoLORvhyx8Sd7tlDKN07HUnRVNtbkFwKzlXzRw
hOhfg55knRZGGHvYJZnDT4IkGOvlGjj58kBd/x45KG3Yj5R2Vj8vt3ou07mcoDqGbLyf17ePJhi4
eMNEzz4YtT+h/FDnqVHCKzvbNVBvzKSCskzw3I7WKNkxY8u6q7yeT8JzznK+GXTXq+1bB4i7YK71
4M/tA0hXVJLRnkiDQD7v40Ej3AIlvn0s83AbaSSWuZv+KnyDFKuBbxvsc77YQLlWatHHUXGUaCCI
mVB/gRmihkdbCnpFS9w+S37bKKU9kO093xcsnDZihfQJtUelpt+0o8ngm/WXMGEWOTHXNDb9kmEP
PrQFLbkNom7NmTDi0mrL+aEs4ERCDYoVX7a07NfdV8aC6cGnMylvswOLnZSh480EMJ6UkQsD0F4h
iMbFGsrkNymRhjdK50XDTbMHzyEV2ijRiSkwvoqY82URlCnxYuiuBIc4U/XS6n22i+CUPBUPwShf
RMLUr+1pk5fi6Z2Y1E785706ijS0l2SSfT0eQGpKdQYOQFjANO1vjbZfczIHsc0Pmr1nmmqC79mS
jFL1g/JiFjGCeEhLzNaBPemIKLpLr0zMBHNPb5Kjht6adRk2zl0H7+bjojKUsYNjEEnXtAEAggfx
iLgCgzkq5jqXKSgEwLQUscA3oDn6blwX7VYIQ4WNHcGeMJE37lZfD4IXSHYFRg/WQy/AkOWRpsAp
px/ek1lCmisUcCMdRhi2lZj/AHoEAhllwXOkakCTR7vouqzObOyn1g5M31m5UgwOUTj45hyRHuaO
BCb3+Nqp4YAYihNnGM1LwzQLv4CJmXZahJHVhUnx3arsenYIlfjjFK5auH3IzkXBmqf0f//rMK2i
VCAysoYXlP4SvQM4HAyoAgq7HCcWVVDn+fsPGGR/AThuSxhzFvE29ipDIFpwbOzeYlImUn6OCdW/
3vwxN1tTUCe3b8QlndeE0rhK4XWnWE8hHwlul1t1mZwEfcBcNejVzxqONfJE9AZpuCCBtGH0bS0K
2Y9v/ExP29Nd6tbJGr6FlW5QSPL9oLYgjwoKSdeHA3T46mYeIQe5baUNephCwgBgOQW9uCnuAR8S
mfdhLi1ce2QV3eVwmCFiAwA+5uv0CbwpkO1gS7grvUqDSHm8VWAxZ2auIrJGFPnQoAoe02un0r2o
szVDQB4cxZ7v369Kvvecl3YIlOxp6segSUxKYc+tIFwYeIy3n4fFzFdYOA3n7WiYlOigJGLPqg9k
BJTMiwNLvG1yVI2wqTDGu2mXEvkUPP0bKEbuuTgqZ1IBEe9MT4MvhbpuA7f5sBqTUR1cX02cWq16
HLw34etWvnFvl1s1KOC/lE2yerjVqf7G4X9+29EEepStnEfUUkfGNyMtvPz1OCfay174Ul6ZJBcj
pp2z3UgaWGZzA1dW88zhb6wCG8hm5V6vCEY11B0KiJXw9VFdvhRD2geItxNDlqw03n9+Z/f/bzc+
F8G2zdDXHw9kqOTcdZrpTcJaaXTzIPlhqnVG54QDCsvW87BuoDrGcTisjlk+k2Q85pjOzt3N3Xbg
cHe7amrirueFJtnjRnGtVfLzcfNrVpqASbffa3WYLUQMTvHSGJQN5pkXkrFM1WULCRZdSqyZ20T+
lV6x7K6xuGGfH3u1uzVOq/8MlKCvP/yh2ivpt2Z0pfln+a5/sK9VrnWuz9As24QOThb/YmxZSKSt
vv+j6zGUAKiJJn04K8EDlwZXXh0YXTjbyFE5xFpFHOhCSSF+nDWTAYmR22ATmM/xwFbJ4StraRfJ
UWP3ksikrCpUhMhUZGSpPyKcHbaHYc8PxbiqCVpnqZvTfW7qbR6Ck5sw9mmbZsR5MVQFrPUFDhRw
hOmVT9C28TEmdwUknUklFI+3MlTS3DFhOIbS0FEAUuPAWXP6DIa0/FAiZbaLkHUWia/srkWj9V2d
VFgcobPnFUjtVMN2aKBHUnd+xBXmjdSc94/TdmSYlXyEFRAI7CXu2poQxDvtLLK/E+nz20jytdhy
9ll5LGBsdihu5ilWHcCvyx0im/1UHFyAgRIDdfT8PtcWnA0jGNGTb+QJ0QB4CZabkGVvERHRFPG+
oyBnAxkt2npDKKfNlktVAprGzczx3Fu6D6W5wvxtCOBz1qDfmLKfIsh44EN0oilOydA0rqWQjMuZ
hit8lomWis6pDfiO247xiiLFUJGaHXpSpTPul2lCqU8twkU7zR9sRXUmrqb6hDrwCJ+gZDfuBwXe
4svmgPkWJEI8FCAO082T3WB4ld9LDOlblDdOIxOdrvE+Wp93rSnN8+v4M/JmvvqCDK4YuU/KW6fh
lS1P+/rI6NWUVHuu6PVY5uTnV3EqHCaZCGbcBQ7nKuU4x2GMeciBVj+3WCe0SYCY0IfCDn7BCGRS
+tyfLAnojDmeiSIfHaQWTY1ON/BR9rDLpsCJ0C+sxEr0FyTB3ocWA6/otmoczLF1reg4tcM007eQ
ktEJgKpXDNLLEIldwM1/BfhabG3y+XxwousMj3dZIcqGniTqLFNe5QB9BkCjPpes2QBNLhMCPlYU
WAN0yCfaNFCGPO5xejnDD8wH2U2QZSOzBWrSue4pxw9VXOwDW5fx1PHDqRGFmFGZ/WI13as27eip
mV90+ftvxbFs9qljwoo62z3lTACipO7kg4ecSrv235MUFXHl4afEoVXkWpgJOOvjMliVJQIuTOmL
H20bAoiOMC39Y0OlrrY/i+SDyaKky2uXnCiRd1ZjSrV8uMdIXtcOyc7/x4hDgwQ36IqqCBssdCTo
BSA9aXQ31KFQIwDcANaenbwIUZ/ovp0+E+j/HLazcFym85bY7Sp3SoCMpSleb2a+uVGit+NFWG6U
sQIWsPjPpqvec2KBbk4InCx6f3ILo58jfw+zVh+7pNWnbbtrB9/uVSCPRfs2t9MHMXLNnkucgWOj
VCQfEkSrTymwkI8Gb3MKnoIeBwjj/AD4BuSQ6RNQoXVCdn8OzeyHaTZqW/NDZ4zhAO6KHPkfKp7Q
NkYMPiaTeEUTNp1i0TXgml1mvIVgaTCQG7gpYy4OoyyBkeOD25WfBGsSzE7G4kzHAzCAE9mpbwc8
CITbrPjhrdBnJ2jzGd9vHuMpDmwl0OB9bjUKtOTX5ubduLgzdddgLSfKoR5kKZg5SZ0H13Wpa8iQ
vwovbm9lvHUi/ReG5fizM8szsCwjPiKUkztakn7SitLwnvdhPb7umgSQr1TrxVdUKIkhACA/vAzY
qbZs3nvsCLNel2A34Cs73uSQAhEVXXk5jldAgLm2y7KVYwgShYCSyPd0oXr4q+Ntsx67HHsZq538
BDUVTu8boaqNIg/kyj7ZIMKgIHkquzdqEuUdpjybicefkAWrXKaP9KHwjy4Ds2qChWMcoZYMwCUj
pjDkmLNfThD3lMqdTHd29qq3s+en3B5bo+Y8O1zlUhpm1u9qGz4Fuusrn6CWy64zNDO67vP3oI4k
cU/kU0Kw/8kAfLVrhj6aKxySfuL8P0i2LNFIeHsm0+ixqOi4YpRe+ZA8TjUDHZUT7OkLpH9nRgr9
Kb8mCGUIPV6vBJXAgA6WtGj5RpIsGumMlFqgWuXIwU9SvbcXVH/MhYoyXesFLWltDDAHwgY8MuT/
5pd12pgs7HjsZKfx0Xf625Q/s/qGiqxxpOAQgvOU4sv8HMclrwH/Fus8pBguNMP0LNhcFwK5ZvZR
b4s/aWjQsxb78Fa7SmMZRpO1UAdWfwaLwPle3fvCnhVottHkIKSU2NJmIDdKIC3S2PIeHdAciotg
ndojZL4Av/xzwk64u7N/yDTC7HkxCMwo5Dvo2d9re+2SyQBO2XBQ/6GxxiC4NOinXeOQtJcTi9yC
xe6eo/+OEcBJRxYZGJuiInZaM16j+G9eRg5IfLfZfyE3Z/6LwYPwY74fZYGgaAA3aSglFJfv8mqe
iz+H0vt2jpEuT95XbAf03+Khca57VMscIzOblWxvyRRwrjB5LeuKo2U73On07e4UEfswo4yDkkse
VoC7wRAWrVVwDojY2DISUc3wDZ2jP/M8E4uwUHgVX3JtFBK5R2/n26k3HsCz4O98a72nQi/tILs8
CLUBGL1vnQ7tGEDVBoC5vcVpmO1rzOKZAdD9ygIphBxilnum/CQbBvEyDsHQvxcA5LhuNLhxZj1w
SmHqLpV3SFKpBxFFTPmgHG/AUkPae3wyWRUl8PjmRiw6Otm16KJdeZlMV7yc1zawr/yBY+EpzuRi
jxldCzp0yVzwpYh/5J5TGdWBSn0v/xJk8uhpfeYRXgsRZsDhEP28LAKvHBb8F43hgFIJGJ5M7DqV
Uawnc6/vndXueI9D05tkkbJnHuCxg1BjpUUUXCV/hnDnd+VocmS5fWeov0yr4fPxZi0rYtSve5rz
qNXHj/IlfvC+VLWFT1je9MduvwICpHOIHOE65eUjpNJYIsjFPLSoWEF/40gBXQ984mVDHQn01CrA
ABxfWzJ5EArN0QF/Z8plXqPhY0vEL9KPtOJAYzToWTdsW0y5rOFD9P460bWI53He5kL3RQkQZoUk
EkV9DWjcEzPCqTWS9AIKIn2zaZHChEqcviwSBQZD8sGVMo6icDI+TOHZ30zVpUv33V+8/gopuwAh
O0mea0nrUxJGBK1MlDUIY+GmfMrsFLEfK37Xfxv3GY7jFu1/NVJWuyOHSpQ833knDmOQGj4JPoPO
gHvBDf0Ss9jDeuFQKzbni+NeRAzFTnaLULGOXc6qTkn/ymObTLpH+d7TaN79bB4ivRLwgbi/LN1D
7wHDDkT0EZnUHL7pScg7pTy6fqtSr6/7pTZOBqvAz9XThxdFR+C++APv0RfceHOw4GHSh+JRepzK
J5L4bdKiSlZihPaej9uTd86iMRLl/AhbzsZFXtC3QNYp9pTux4zBMefeKmvMgRRoUL8wu9C91rjD
f+DxJvtcLIHwy2rnX0Vp6M6uvvRkctbVpqaxuG2sL7pxm3EArJl3NjPumqZH80exv0Vy9XkX5sg1
KH6i3rmtvnn8h82xxUAw1f7Z05dezfqorvB6p2RfFvK0KBtUfTHLnyT4wSoFE+d9/ZZGCI/QImno
mnjYfmuDp+d0rDjESt+sA/W1zkzqAhNY1CYlDAb/C0xZC7wU1iRG8B3m0YtpXKYREF0+HYmdZQi9
JJ6U17SBGuyuA0baH01BnB9V+2t/jNYH3XflA/N3KjJm+Eouyld0fIz2BUmu08Yp4J0NNpb6nBZX
nY44vBZiaZ39hqiKG4cZ/NimswrM6X2gymW+2kFGR5nbJ0OI4EH+XUHEHuH/1SqvpheYch/aQEiJ
kx+s+w0lZo5w1g4jlH05G0sm1mM9o3I5LTngwS+TYPNH20tLswGwWGyPLBgp1UdWCoeJQCUFewtI
oyTvCc1fTqJoP1oDO94e+DC/b+vwOFUOUo10/QKLLLbaKFAihktJh2CBKZIuHNijUux12dN3rCsl
efmbyo8Xus8/iUSZs8XZnGck4N+Mid0MxhAhaEa4HdjPLp8HrdCWBLo1bFGoVwOno0aUwEP9GkyP
J2hekNHXBC5XTGFhfXvG0YNKE9AYpQxM1gw5fzGU4RZn767FZHZ7wL+tA/B4hzkB5dtvcMTYTWnN
F//29lInHDRX1yyozROwVr1d7PqCXr5C7LPPZk1loNTRt3bhc+gbHwl8vXBy4z0G1S+2gyIDbuOG
RxsuM6TVFzXksGIYr05UqrjUX6GZfovT3oxNJqjF5f4/18LN/cHKDkX9eETTv84q7f9j57HRIaLO
FegNl1Enb0fKXyurQiR6vS/+akYqTZBoSceOh4Bqgjn45GKxGGCkcz4f2TAUOY22r2UQ56new2xz
U861Ay1V3DQZftuDvV0VPYMjn3SnSKQnLFYgveGj48P4FgrfOav4hkHw9cQNH+2IAm/l+irfueuj
IkR0Vtk/CxMIxGOINhTvknwe79d2Vl+VwQbnlTS/BFDc8CXdpXFkPSHFT2J3Ezk9qNyqj3wGKU43
c2kMGK4vmfnruuqckBcZdhoAAt7XbAHG+Y/wt2GlC0Fu+AgcJBmjcbgIju0eA4W3imet05Hh4fXH
/l8Ze44dK6IP1AYritbWjIGn06dVzavoPSISPVZ6XJxuh3Dq20rjXijd8jWsfLN/Oxc6TqLSAIdp
Kom+WrDvQ5YKolqC0PPFQlJLeHdZ9vfhfVEBZti/VAFWKYZfwFigv0S2Kexq77oKAgCf9/ZXOHI4
wZdiOWdqAaPvbM5fCI/iSPUhTIpYE5UH7bZkvmayw54V3AlVP7rFgOcHoqq6r0FVmimGtjEv+G0H
55qo9cXko51CenKP9bcle296bS6qMNe0RfZ+cpxdDL+YgUSrvYLOWBFuuVS1Esq9btI2H/3+37Ns
oQflGsHFTHvpIHbdIyGck6rJ90LShSv2UeXGekUZXax5G4oD1AYRPqKhDVOsvYVTwkBYFFylU4bm
JDGNPLhZlk5uMmiLRdV6ZpviEB+C+EIaygjIcmuEhmm5Sx/+nr49dcUKXNjShtE5F5VhzcvQrnKQ
BpNQYvxQgz7Lq3vZhGP2CUE0MzGbQZl7u3Jkk5ywKlbwaoNLNqfQ+pe70WG9pk5J9qHHpeaWwwo5
wIuePRZQoRB38+RqjOYsFCG5v/beYywEg22n65VPyBdzwsAHwMXzks5Be8WWbxKLw8BfiA36Iek+
tHvvbDdQkdxOdR/hubYzaiSyv3qG90NOH5QPjxW7igXC/hZvzh4Maxby1YmtGJUrqvfoEIIhvuty
4g3noAULAU0iCxEFJ+iq/pvv4IfxcUS8Ve2ib6qXohP/PPDnY59U6ITKVUoMKFMPnobRMFZvcLbP
c3xqdHWWA2mPNNQg9JGNsKjLg1ia7/R/BET9bx/7Zz9pJvxEgyE7vUbtWhf9n4vE66j+df9cvEZn
II9WY2sh4fKydkdqpOcMh7e14AlkRfw4y5gRDTsgUIhcCn5RNgNTpivAzRnvbnshYqJHiOIrRZ/T
W/d8K1/UrqtPT5zC8k026+g5hAzpkrANyxKvNd5cz5FfJoK1zts89gaAigscXyQ2mw/KOKtp4dcX
q4ttCtVM4ALNdbPfM8siMZnOgL0D8NCC45WDKrAxP33vtPFOZgPHXRY5ui7s4AcrwziYayFzRvIA
3loZa03k6XuPclbgPDz9LAsSZDp07vP0onLy596ANiEILL7KG4gUlhZzN9H3LcrP10vtx75HkGcT
bkc5ROqKBCkxyONIzjh8OxuBH2ilrPmWxAXnKb4rA4YJFtl9Y41IlcRnjveQY7deaNxGO34HesF7
ZbRHl6nvGKPveUVxzoBfYzYSCrNXDoaHLpQPlv64a6hTc79YhSNnAKnXc5ZYwgUgba00YCvDMWmn
M+9lOlJh0ysqW7/CauMi6kPy4jAVbuzpIvQirmthvsd/l42ifujms5Y4IHKw0cI+ApZaFrPrf1c+
hWSDuGlXK6MInqodSGmL/n/k2VFQXNBEtzJ1H22mdux0bScAwiYTliwFbuE800W47fM869JPn1/c
+UKMUuAVL4RHfI3l6VUlHHmWTPSUFiPh2buFU7a/twHDeb5Jzy8/kJgTGNPVJilxJrhb5LjxiZ45
f5FzVkmhkgllJRI14Cjm34GgGh4z4hswFCbJTVxflB8eOg2s+RGI6JeOYm/RpTBH9qRad3oO6Gtr
uHZVQU1Pc/2AqE+f2BJsZKSuUTxOV9IPQ7zjIXKoBy2lD9qVWWnzr6cyBVDG8O22HA32t0DJi+hh
bKFQom7Rooa1UxAlwJbJ5GcmESv197VlI3E5Nb09M6ReGRTiJTtFXRR3hHDxb9zJTjcLiFxSbqA/
Jam8g/ClVOGctnMmz9tQKYVLdydYLRGVdoYKtNPgf3WY7xju5WGTKzpjgunsCpsdWKMZbbgnrauy
W3OIIsP2ZHMcAPg/BKpXXpZ+JAltIRsWcJ3K72vQ6QJuNKRSXUOKOrMyrYSTdMy4ydF2uaSpKij1
JyXbOC14Bruk7wGV/ELoT7bQVKZlemoRpc/AUXJjjyu8RrfFL/ouvsXv29sYxBSSu4oo8zOY5QX2
jQ+q/qO10GtszELhRf+pTYprSfzimcK1W2iWLfYNkZZ6W8GfjYxPUYJ7Y+tZ/aEPotH+aAYG1q+d
T7sCtTNRL7YEw9RQWSPVbumir4+OAZ+Gi6vs0XgnRrpHXQuZ80gG3nFvJ3EwaDszY3K+xBrsrCW9
g6Q3IGat7S0u/jJEv3ScX3NIFSWROlQyBC1Bk8e/ix6HE7VQWisxyiCqPA8RfemwxIiA7Mqb7CW9
6Z3SNuMJ9RoTCQ9+9L23/KwadJASlTdcxvSVRQJyxGT0I5gAGqbqYYRqV3qhLmpYMTyrlmezagcV
tcyoVd6Ii314jm41R5zTEF5YqLI3SXej2BDSAXYmjW5C+wMLmqSdXsnY5Wkbp59Q6mDQPGORtTu0
PqUkpMVH2h653iczGFxezzypkWTwz2LMP26oHflY/7ChhXoxscudHNcFA3r2+ArnlcXdPHg2KbbQ
3l+0KGMFfZqKzQA2H298GuUgpYwGX76b8k2aCanwqbQwOlF45k13WD9/xMjcdUreEiaA6pqt/vg5
1MreDURGmKl1Bb5GqkSPmx/B7738rXZILhFnD4kguPCTXYRH6cbPFkev8a9q+ZVF2z872elxI+g3
22wLPciS8QpDIm5nSrxF7/E2nQE0qwfnO+7lNVRDQtUh46xCuNoYYfhgxPQsmiT0tyyND7dbSlco
pdf8sTBWvEMUY1DBFxKk8BZaeQWGE83wLCTRVBlh5zdk6MCPNlP4fT1V71jDku0CvNHlpw5fWGEk
09wCVNaCrGYtmXF7qsy+Ru/f1uI5mW/jVlWvtI5WT7VRg1NpRWnqUDM9DBKcTVRmoMaFgInJvgfQ
lKN5WN+md2N51Pvwddf5dLzlNT5ffT/+akqLQ+M9s4r1FflYUBgJdOXMTW1y9shdHpKXAljTsg4W
oi9cQIHR842K30p46T1Or8G5e8Xiv+cW9gU07bbQClInM7ejnCz8gnYBt0eT6PiaqaastCvSbyrt
fe3v+lRp8yJvUsUutzsmtFph/zFta8q0oIoXqit5fUJvIHpljamqJTgw3OAxLhNMWoT95cU9INyh
C7Ir5Vltwa+HOOlj4623NrgPYFPlO3ODQ9268a+xFrh5NSF45XNHpy0Shi2RDZJ4LRli7Lfk8c3A
pvKbQxpSvTjWFUsdsnLaYXY20EraaWd6oaSc7jfC8Hd9n7HRucwMD38aOnTpuvXHH4BuXAByRfwy
r+jEgWEjDXuW6KbcvAaA4SpP7kEsSjGtqfccv0Q/GYaqrxIuFqUMh6nKKuFlQm0GpLRFevHRFU5v
pqz1tmd4Rmvbz4wov8iHPEshGghCULi2irSGKOnhZO3cNMf2GzfduGa39bVkVIYTIBg+ynRJKGxT
WwyFLAvx/Qrxv/+ZXbpvtS+DNL/qAfiIGvjHbzfI5QS4dZt3wCMBn6UR8kg+d4JN4aGFes+i/TIt
9Es0MX27jhO2FeZ2HjcW60qeZFNEudDj6aTo2EiDDoXfzGdAw5245DrmPAC2eLBBoh5fRfZECVoI
OtmVn+LgCLsU/Nr5/op9PhYjDr8WZvTRcW6Dx/wkAQ8UfFEIVC10lTe6JbRzzNRgCwiNTfQmpMvn
L/s3IROtMn4+oSA7WZwVg5sTUT0DaebpB0TlNYmG3nuK0PNiscq1utKwWgHByjukbo4vPMPyzS7T
QeKYsMuk7N99pYp6ymG+3wSjWGq3PiUcnBzLH3QcZSzY/snGzHP4VyeO0/0NcEmASBFQWC4BTOZy
zMeMD06WEIwkpHST8TiD/m8YIRdid+WWEwXiWb/FG6IKZgJqOmXUhpBM9iMZGeKfZHv5lvcyol7A
je/vwLa9nLhUVSx/Tjsa3qVh4H19zjU0IP6VYCPimTaijREOQuP4hlkKblu0ikXMudm0fh1M9Vyc
9+iUCt19cT2Cibq38KySiYUAkBoVIRJwc2gEkHU/nqwEySabTNH0h8JtuGyaAY8ydEBeYPh3n313
1cK9kqhM56rkhVH3VlF2mf6RvKWz73H8m1AMLRtcwZHXNxStd74jjTM/sm6UTQTy8ltfcg88zgFO
4+4sLR+asM2lG7CwW+//QS6SNk8E/IsEXaNdDkJOBBTqoKPPrx52ZS9JlzGaFIOXAsuYVMgv5git
U95D6PsqieuDGrqcnDpVFsny9p7HJwAhuseqlgR/Vh8H7XdvkeE5L0nLgF3U9pxevHbyu8zTHyvr
Tr2Mpmu+esScs6g4eFpS+We680onp2QPrOS0lCI4/8ZtRZz6ok8sMz24UV37wTXlaP9yGQGup89X
+Ey+SulxlHMIzVtZEG2w/E8uvJUldjEcjcLd3W18B4meFGN3Yo69Qo9qU7cUeMKUAeZG5Vm/7p1o
TUbk//jtJQug0+gOUKkf4OHdCr0M59qs7vAOxt9piGcF944Jncst2rItWWU1c18VWSU3rPf5KZH5
6w8tuEjwuXVPFBNsgwwyLiURMG93p36+eYPKBwfngIRgmuuwMjSUvKYrW6gtQADiTxx8pQdhTiki
i3QJYVuOXLXdoLha50cLDynNaJUPZHj3pQMqcnhKdIgVyJotxl/t4KV9O1+uTfCgaIQsC3Rif1kN
ae8agpb0LXhtv8q5WaaN5Ejg65Lge6C9c1Be/lteTsXPBbZYC/pMbAlVTBDS+woNeR+GB6z4PqPH
TDdXJ3lc2SRMnjBnuxrSsFJKPL2oLk8uaims+2UoywD9gTnaowoto6Gl2m2aokiq1x4tZ7s/zo81
FR/ruEyZYlhVk1VcdYLLrND2DWQcMQ10cf+mAcC5J5LzQMyp/R+N5EFsvqINPYs5CEhLRtwH4yEG
5WtwN2FAZ6+vdp7zh3LPxjo2RvNOny0ptqt6aRYxD+2CaBvvx+iGMfyH9/TB8gntgHmoVvDw3ita
ny3dB5sIDtSXHDysJVHfUt2gr7hhGoxQeA5qiqxqS+d84NahOcCDKQmmZhWesDqhqmH7w2Jf0HiI
ZZkv2GS0w6GBM1RcMQSBHCBr40PzzE4p23X0u9xTeDu1VZ3Kh3rb2MO48XickLOTvWemmJj40oZL
wYx1nERAr9rZUfJuMO0QyhGnwsYfAhYTRBZMWdX2b9fAXZsVhmv3QryZAVQgP+RKq/y8veOZQzEC
hWqWbcqJYhW0netu448pRpvyijou6vIYZ5N5/ppGgfuTcPIrxx8chSmDhZShtFyKQNzOQ4F4P+TR
nmuZtI2QHzbdVsctYnBxcbYZ3st3CzmbnICDy7LPZj2+6sDbm6UEKRpQzkOkw3iGw63IJnCeQBIL
s50Vw8fSYZNqSethkr5XS8Jl7eXmXWIUrGSO/pwEGI2QvURDgLrd1fz8aF0PNPWYqsx/KxsWE45M
a51cnN1drG1OxnxBUVxkWO3tTCk1E+hdVdKVi/Jf4PDFrNjq21JkJVFPqpM0wFugXgCmJq2EJaGY
bXHYlabDA55pOts+q5OZc7uoBVH0QarZMa7FV7A/f0kGMgGXESG39cVO69HpFUWrAb3IGB5etrtf
4LOyB1EJAOSPpBfWmoUU9PMXmlH021UrmDUQL2HZ/X1f9OkKbU01PDdGsKTxLC+IY+wPe4m0StnC
BU2Fza8r/TBPryqEsRAVVqPw2helFkIGvWwNghKKcmToZrqaNaGxhv7cObkds+un4kcsOAkSSTpC
ipSCQ1ueKcSjxvO1UMjI/CYT77QbOTfcqlbR7HRUocVlakcRQAhLlXKbJpDpqiwsOQjPehfQlM4G
sBWxLV1YrXs4KkDu1xnP0Zt85bJGqvuP4/z8T15BCQHz158JlB4c26rUrCIM0568/TFgoYAxEtbX
djA5vrH29u6I1xMUk8KIgbMEEVPgz8v5JtWYuBrvtsoHc/VbQedDxkBHrhlK8XlJf/rA4oRyIG1S
r/WJ09ElUd0f/g4u/LGkc4zXsm5Eyzk/dODa1zFBAlH8CC7Z6dO6hzMBSvZWgN8JgL5j6J53exjj
h1sC0ZfhhhjcmdmPS69vDD9SMfY0ZxNrqRq4dNOJKKm8VAbxzvMb2fDEAEyWDzjf4+jNApPf6egc
8eXb1EMD/lOel4/opZtlXoL0F/g8a06RsBRknfAlLKhN9EcB+pNj+9hGlwVSQyiW2fgs1ffj3OAq
eCrBVMq3XAESW+Mal+TO8EHDdpMpC/OKCE3noxoNsMVltFS8y3XXSNvFHlvVP1ySsEnaWHmf3ZZY
imDcYN5Df2oytrOMo1Mk9+l0Sp2mR2YhcBpT7/XTv4z4HLQakVMvMHLXnhlL3YBzeLaxOoYpwXtK
QN9d8PnC0mRZBB5oa6AYRhVmPmrdCagpNk+/IlsexvD8VXuRRTM1nLQcADoTxg6qJf2nKGazT3Bn
tCdkTyBCK2aE0YBhf3RGidNbn9acUtCtpkhphbSrCvQo1jnRjq5FTeBdgVQWLeyhkvYKwksJVFKy
lj/QX3cTSvtrDpSD4NZeKHpJvnISIbIUa+rMrcDdp8XvlydUjjQFmjHmbIbXxo99OkmEnI2hJGU2
SWoF3EQG1gAOsg4w2l8Kxe/KtX0tg4zj7RsErxc1EMMoiibg9wRKT7TO/3me1XK7d7N3o6r2BAo3
c6JePoiMhlEdHz/bxPPajLb1XvXXxL+xrbR8FdMkIhUnKc81x5wMT7r4OuQ82qFojw7Z8PIMrvhl
KxksRpxeC3rGu0tXvhF2f+FqbulPdCBonra0zpK03CrI9qLi1p4k55qSsqQ0n9tTolH92Em+03QI
u053S0d17tfOaGmiPHsloBP9iizdEBfY7QntKXRBR/cRiDDTBAac50B/mbLFUNH5mSFe1WDwKYkm
92szEKwwjhHGplb0m+0BJ+A3+uguWYUkgfe2nw64U2/tl0UoRg5KVLw4qTDgXkKgEY6JxkzKpUp3
W8tihT/09oZVVYwunOagApvukA4X27EN6A31Xcecsl9O+vFxIeSQaGgNlzytL5CYKMObkecEojqH
tGnpXKfAlALSOkrW+t+mISJjEqz8MA/Fd0+ptifGTH9x6yNWrCCSE9pLL/6PryPu7JCHbcU/c1WJ
eXNaYEGsxmyCzen4VROuKiUWVGdiL7hcK+chExYkCLqeVI7YtDlQatGezIrpcjn5mM42LgWp3Uy4
OdfyS7fP3YYwXW9PhtRaDvYnFfmoY+97o+AE+Jy1F0qr32JixUZLf1gP7GwbFXIXfDrh18KSaeAc
brHWKOe5srqqX40ZuFtOX6LqwfTPE8OGts+RHUrZhyIXoxbugPX4qhcsD6OXHh7dAsMIVqZXtyXs
mxvMQS4Ns8ah4RcFe14OouXjxLr8CvlCH+DgiXehiOxUWZ8cCIjMeweRSZO6ozJvocnPudruGxhM
yvEdVQtAxPRT3n9wJeOIzpVSTRD0q0G2tbop511Nm+8KzVvj8Zd7/1teXzWkOwYXfwu/AXCcNwW+
i5dQVi8iY3BsdQUmZoiio68velr2mIadV2jyj2U7X14tvysAVBpE8kIeUPTqNQmTSJedqhQRniTO
dbNLaA9tz85G1qthN8UifZ2DuQs+w9AwqZrfA9vTzX4UPfYXRXSijP5l5jSvn5QecqRGevgXcV96
XdfDS8EkS6zGLzPIbWIyrVmAN5tTfc4+cSeib+nnp8a6vimA6sfpc2QlXDUPze5+uSJVMyP8O0rP
WX31EwgYqmZpAXI0tO/FnzE3RHu6yN0odgaNdCgpkSE5KkIR7pEQJIHzZMaB39HJ4wY+fh205WbZ
5YlaSE8jJHB0bqR5atEFcmmcxeH9hWf7sIl84nqnY+YDol54g3NxOaFhawddF0K50wtOm+jCiL81
HmANJIAo3LYBGwdIzPkfnnrcMbUlJOztwEoaLejRM70jZQtxsClqTANhP4JwMaDnkoskg+iPcG0q
fPnEv8D7cMHTvuX9RrmDXA6bf5jODLmqDww6BZbA8sJFCyVH8ZRuhDA4qKnRzCVjj0XNWRsHsU65
ANl+Atb7+6ie99j7kll0ahp28lLsXysDtvW8RjoI30H+EFstxSJrnCxZdo5HuGxnF7THybc8C6Z2
tB8dL7Q86v3Atp0FsZVRHPKRmq/bE+dD3VoGWfswpirbcNBBCW7s6iIR6HlY0DGhv2utk9yNDUwX
Vzu1F7EptfIJwGZtSLcOrXfhRE9xOLf6vV2IDySgSzcf44t9SV33P0ILC+PPpxZ0HAZAczORJuDl
1BjCzScI0nCOdIrvf0Sc6H+Eyad/GHEM9/iievnGwR0+O4I5+R1jJJiRBc+KC99tG42WUWMGESzE
yuzTvgA2F67Nv4cPEz6ucqo4B3QZHsmuqM2JXAgUj7Wvql0TTIjADyj6fBlUXj1YD1xvjLpZbO0v
3v7uSiYspL1uSO31Ubj988Jg6hN/djNwQHIMknqJeDMJSuohlNUvpB2DKcyadYETD5ZrsKGzo4wm
juEFq0hOry3HlGLabHv6498fIglgpbCwe0gAzwDcSVUjhudFgMsgPsKG54RHD/rOhkVgexjM5ioL
3pTgiOUyKRLtOyvV5KaF4KK4BkLxl344z+STCcwTYa7iSHYifJsTQASxjjhX7m6jylaYzpuB2xzW
UIq4dOcMOWnXR4fstlQtdBoZVkI4T/Gpn5iOXOoqVt0LydQb29PM8YWjEjkDp3hbAgywVEGEj4X1
ilPLRREFaaIl0OcijBzgb0Xk0UnkqP4mXXBBmJgRXSylYx8Ks1D4J+hbOHlhBCLaf2Zd5Oquo1qx
E8/EOmFnELtvxGWHLaDtodEV7WGSjN3O1RvobB3nyhqPM1pQTAOrn+ZKyystXcW4cSdn1yrJ/RGF
H2SucWxzFGGwpdhdbd9hVPbKPtZHTACdlNed0lBqBOrWMfPKKa/WpBzJSCXDwWGxSsNy9a27bCSk
L16IsfFKsr5Jz5jpPfUKOtLdnBrJOdVUwvbd0/1vh0JP7hHn8tgb0ehrcEECnTU5pQsWGLrho7lG
daOPzAjQvDPgb7qC2n+JMvso9XvT1U/9Vl38DIeqwtiGpTLqQJRZBTXuZX/JCYeUsHtTK9AuZoZV
aFLCUcr83K9zrXw/nKCUt+zqJesfd7XZ/zUb9n9GXnU83iG1digndonL2M8WFjbkCYSL7i11ZTks
IWVnEIvD37ou0i6F19nck1HdFtut127bixn0itOvcR/B4tnL1pAWWDoVZ019tf2v/AyaDClrdE9t
+2L55JlbT9hVbuqG5IFrQJwuh1ai9EgAD/LuRvBVR18ij0h3OzlhC72iRgpgF9nlTmQg2RpXlWvK
nSIv16aOUj++Z/LGNtg70TWealIthA0GpjbPanWeX0pC352nRu9CkTW50XCHPzdOFTTbaPeVwW9W
SHT+wv7YKkIOquIsM+j8ZXii/h+8MBARMzKhja3fswZgz6ZmY6KG2UmIr9BIa5egOkadolnmSHsE
SZaJy8LmF2CYIs7sDybehcGvLU8tsA07hydOBdKKS+S407BeFkLR1GgcbgD9+UEGAvWqj6XQ5N+8
H7TJCIN/5DM+sU75a8E6jVxeh+bMx7NwEnP8kV9sap7FUivGOnm/q0id5HIkGzPXkofD8b6fGqPs
qsnorLvw0hSlEWrFtOuT2I+wnfuGwMNLfJpNrpC1ZSgca/ZvSislB1RSJtjjKGEPsgld3S3QHgsx
HiJcOvcbkoBCQKy08GA7zXs8Cb4p4DCMlkOEp9nWGEH98bZzHugMG0SxpS5DaR6dhYqAvtRt+VNd
6asd7V6uNwSmlqp3Go1wPsBKChAwA38pN2Z2QSlAyK+orQRZNVwWuf4Crv8OROmsbed3L8pOGC60
btQJzS1htqwsNBUItZTP8Q6h6pnrbPaZX92ZPZWxdHofRt0IkIYbLhreW1eOnSTpv/n3IqkDFlde
4OMwRSkwHR6XZ0tjGeK2Ac4E9FF60/pFnntdqea3Alm1i303o7WpaD6Qpz6ST7VnQ/GzOBaZ40uX
JwwG0U8r2G+URvWQBcGI239TmNMW2l8gEmDLtnl/9AdjD01JdXno8ju1aBlp465jZOhfkEOEVVj1
MXyTfWOtToKcUKbTzZVzV4gXIaJnsCa2AtUWxMseYyVDXWDUsEAPhy0GpdSvsVt+DOC+gZ9LiIGO
VJUdwPaijOcJeh7y/reNLgVA4SvVPrFMwd5zJkLeb4mvxe0XxX3gep+5QseffmHsOslRSqX2Lrhl
oGl4EZbxTDIgLWxS13BRVOeMkjAwS1zG+WhU98OgyrQnVHK3SdKsm1fKz8lPWfm1ku8nEouzJEDu
sye0sOkHdiQR1RRViMKqvaSaBsb6vDcq0BOzpLK/r+hnjvGLEC7oGpNaPFiWRKIClQMiGr30G7lN
uZIz+j5hrEqFV/+r7y1ojSbJ8xt93bLF5Gi2nIQ2JmfYHU+hquXOYwnLxcE99EEm8ypNAMCFvia9
HwAt5WZqPihrZjil+LhUP/HH2r4dTyALPm91mwX9xI4yrR95d5N7mGq/0TOoOSXVFah6+utBovUY
TBD2Fcrz/abaRTYHNkb+AKziF/SES3oUszZblxiSwYVGkqTBWohlAgnLZEjulMII2sLbRahiWo1d
ZkSi6LMmaw9TT16s5A2SZ1wM7y4eMJFtRgUdcxrBEMEfSgke4KsN28nQs8J/CA5nf+FqwhHiAE/Z
UxFzjyAXliYpH0OzDlYktxc8c53gH8wMSuyBISCDmnG5DlT92hLcQ6ibzHAXSp7oxtwxOr/bTV8x
Do7hloyfUWBvqQAywFsGFPXg1MQVFrB5SGYBD5uNr9TMy9Zl2sexuOXCQtswpep5t1RxjCizpApV
4HFIkQYOX4P3NkIi95fF7pH+Z62xtb8Cbu6+Y0aFvwvWfKnbpb6JDY5Hl27VlBL1Ir6Ux50lZYWp
14tJlsyciYtdXpBCsegTcNa3JtRbvSEbpBJW/Sj8yUB3u7F+qJ8tLhlaePydYIz9GBHsAuGo3+od
J+ypH1EOy809wyl0knR8YQS4mxJ0PNS1jlI8Fk+NnEE+ztE/7x/fxUFF08r7P/bCn00Ytq+500Ph
xxVt4FZS0wrVnhBw7zbhnVv+uXGz4LqY1z1mPKuxiDnAZJAdlVgFdR1xJ+d1q25zQtKJ32+way8z
bu00w4gXMXoGzIHXcyu4U9+X/16p1G6fux+su7pp05P2j5d4a32S5/uQnR19vu4esPXw34i/b0er
KEnj2/raNDiUqoOoddd6hoWzMlQ9iu/GBsGP/vgcKOPi5B5QM2UrJE/QLglnt7430X++3HF5Dp9i
3giJsoca0d2+HnlS+dRJeRwZiiqdppIgsxHpwrhm7aGXjwFFsmQNd26V1BCwYvkZmPeL5rzFpzXN
A/HBQUwjtnsL9dwqNS9ATHBMBaz3ZeN0dKxfL+Uv6zG8CVxuzdECV4UdBDpan2149rjY2Undlt2Z
d1jj0RYP/f8JohlPVah4e6Jo3oMKt2IzS2P1tUNUGqhOem768Xr33thyHnbS0FAiTDl9no9OY5ec
fXjC5JEnOB7x69Ovld+vdLpVrv523tIGJeqgC7n0iwhlend7n1xai8Gd59ZRopM+gn5d2T978554
df7gczMvVfw/IKylBzfdAlN3aMCwD7a1HsNwzMNsCRjs8HEYgvUzGZSeFGllw2ayY8h0jd6xpJLp
+7S6+pICKc7XJF12yxj73jdn4/bTGIQcD+72gLzXU+KxKUVF0C6bFs4Y6Rri2se+p7IZaJoeZ9Nu
aJYyHGXeGuwp/x/yI2SeZmo++aG/TLuO49wTRrYSP8rcBVxo5wVxvC7pSoox4wHv2sTDE49vSq9b
k6Jlkd3dcjw+OA14D/qQNHq+aTu2xxCp10Nby5p3j1cSGU9jUSyCboQons9aNdQfTz8/sfv2Xgmn
vrvqNx8G3GF9vvljxtsuTE1k5bpQcX53p9WP1f3GHLwXtk9XsdlLW0va7NEU1mGBHjUw1vAPnnLL
5d4vEulyFkl4k5sXpThXctys3Cd17KiGC0+dF3TV5TpAPuHCUkMatmrVw1GuBigLV67LGoVS6C0i
mH4X4VBBwp4sB7qbCY93j9FQmNM8CwaFiVEsXcwf8fYi1jKK7q6kRR0gUQf8On6EmSU1xzXAGpkU
246L8QTPjwhSIkYG+SXsSW3sr2W8HaeiDVIJLmE5nTn3ci93Dxf5r0C+fGnJQD8v9itUTAoaIVvU
hvCpGO8UZqU4m1Zj0ZTCRWu3sp2oWBthV7B+J2gj2H3o61m6XIOuNN4Tm8+X31K9E4mQ2rDHvOBF
hzmW52jEo+uP1+qw35o5Rr6YKVZ9EOfYlo7CqekGccrqPGwy0ZxyW3DTouv1DZjNF8sg73+lTynU
OAL5n9Oj/NYE+7toXKs7SRLCfYt3N0G0qfr526fQW7MYSSlQWy5ur83W79R0Mx6M5H+Td11v/2jA
Wr16MfY5hcWbskpF3Ad8zGOpUOFOavE2JsfRHvyjs4MjtlDWhgcNVsfxJBVCaIJFnTZykrBql6PO
4R6vlC4VDTe6YoIxn0an+fl7N2xsXgq8dDMXU78ynUp0wXpzgUEaqElmePnJtRXj7xLMeYvHCALK
BXpJV7W0T/C/S7hw4g3rQv6CBU4qMOExVroJkQ/zNHxPT2Q22RpGWa+2o+ZJm/6njUSO6OF+T5SJ
gE4vYSwlQoEG/VQuYBdAxqjRBHsuxxycaCVlDgaySrJbpZ7oLbDv58n8pgDVIciOqC8OalnzuPlu
NFRkJFIaL3fJgPuK0T7OY7XuzVfBcRcTMr9n8dloGyDdUZJCLo6X1UtDSU15gsr+ok6GAVon4QZq
qBGKE1ERMrDqUpU5yTbvrsVpFGl1JLrSNtMhptZ7/rCMGNB2VqcZ49cvHP1eF2n7phZ+YPKqlJTo
OUZzXMXxCzfHyswwv6lbF+weFlWMt77r0hWUO8et9+W7fgTlTx1hI1i6rv8J7qN++4VGCRTurYlw
zcauyaFfryakjrT5VnxUh8MVHo0dM6Y+9FrUwMzp60+rJk2f0JGAqk5oXCyAJOUbKj8BlB6FUBNv
VhOqmC0fjuK6t81Hg5HhmzEdUvZYbCqwuRZpoLZSFQtIsrs9uqWJ7NacslshhRC8yOWpa8mCPGMV
675/69WoAPfQKQyGmtEjLm4YRMySQTnVpfqS2TOxCZGJm3cSu6utETTZW91BnamAAW3bO41AXW1N
+OQYO6lT0YgORDXBxMaywUSGlnIq4EGEDPDfqgJm+U/7STDIy0HIFeThHQ29mFNv+oJXTa8EYHka
4tveAgustXBfyOo/uDibOkG93ce2L3W9iY1tbXaY8iWRCzwbYn5t0GPRbYMmjkU0mxpBWxJ0FrSP
fdT3K8oqR4gOYzBeUIMVOvZHrWPif2tn0V6OWNAhgH4A5umnxqUiOMvMsnUmdsTUfX81xynHaL+m
OpnVQUXUyqbXFeMRmjIXWulWhtO5UT951LCVdBFNneOT7EEtketB1s6uS+6QoMiAlEreZHtcxVQo
9H3lx/I7PH/LEKjigPEd0ybonGi4slbAsA38IQsXb+D6EGdi8agFS8mjL+DcCKZFFFV4s4KmsrQN
9suRVc9dZNhm7Iwy9oZXbEYFWorENrBHfWvwdgmDfQAaP5IEP5NlWHczyyn4LbZCSFdgNODRCGY7
tqHnZTApj2rV5A5wZOvzp8kioPIGtdb1YSR3SHWxnb/WWhO62aaNqWJTwQywDLOVv77d3FWVoq9n
1dTGLW3gs1zLhb1DjIuDDDSnQnZ/eK4xSiJ1vwmqg0kEiQedNEhXOzbFoB/ff1fK+IFlUPdmIutR
glON3G9XYcAXteb86Y2sG7GmLwheLsOLyVkeVPzxpyj3gtLqMJ15mL3kRnTH18g1aC3d6wjpHpZ1
DlfeKAMOAwsYqp1v6cafzmRYuLsTsA2M8zsFFm0JQzi/Md5OngKZMGYDWMaKvldiVHGcORLAtG69
44a8CPRmSQuOp1mcCXcl4xVScEc2Y2/ouvw8pPKLq/A4W9NOtWqJ+JgDgdWLdn5/vitRTVDAziKL
+0TGCO/4xA9bHQ95Ab4Qig4sSqdBmPjwst2cAxpULDk3mvTDJdyomfmQMxh+9/SCtk7KW9J90Wt5
nmmjk6viwTMrlw1OIeJ8T1SwKZnpDnvEUy7QXPBlnfdVmE/R8JjcR2Z8R/HrRWNmmEnBeh1S8BTk
2HM7BzLpVt/OKol4FbK76xv7rPciRnvxWzIDeO/zFuSFResEcftZ8L6y9hdvuol6WTrdpKZz670b
bUrkOeSPurCEqQY2cjKgRt3rNQKME+eDMkMffEu7hgdCfVRCNW+sqK98eDkl4NK1ijFNb1xEU3em
FIBtvcU7msQ2JzRpSv9egVL57omjfGBx90ruE3zfYXMPb8t9T17PmW8Ls1U2E9V/2lF69t5qTj6R
5gEln0/GTHlE28ugWMhOvY9sEL1JVaL5R7XcJ0kTMute59a5dGMcGt+rWl2S6ElwOAyaPSoUQXpy
EBua6xna4U9BdIrYHAOHw299zv2a70FGRBvHQJ9F6KKStvtOUqUNxPAq7Ypvv4GC4218MlAavtMM
iGmiOKaAb/0tWgvzFm46m6QIJYxHQj2dUvooNKaP5y1qJie5YoCuKJyfU10HbVla2StINRRNZHqm
PWNGVv47MlzjhaO+J8XcL2JKTN2q6mL0pN4TXJOGfZBMInhjzyNUlpvLTVZ9E1d/+UrQqHGTZMrR
8zO25qJhzdXJFpaPgoyfaA6y/IAZWRLxYS44dLX2p2P9VIFQRITAuc0NOdRZzjt2g5/DcwtLkj1F
vPanie7TvQsX6/Lpc0vHYptSmED6NU5SEqOj3sEmlrj3cSJirQpfeWVrEfMaH7vs+YTEXUx1iCdr
wNofb/WjNrQgC3drPsP9TeaGTAnRORgIgslMSyghUWycCszd4EPs6Zq66K915i6EV5biRqwxRCW7
MOtTKnpl649BhBI9DS4ktrt/PACaXiE3GouySaBFnlz1P01ib5TgKOQRqA3ngF+wzZDGGvyOES3x
jKcn6566dVTTUNjgYmKPDIzQS59DYpmheNH+JY/25cscS5humIGcxmpKTz9HmRPzrEelCvSZhuYK
s3B39C+1hihXn2U5CKO2+B/Y+pCSvayGft+/04ouJwyFtX+2f+5NmZ7C+gBqBzKknq9cliVUkOBs
0e8snIRy/jih4248xu+SoVww46sDDR49lxSywD8MlMC4JKBVLE5xNlFm50hYy4PKwekV2kNRtPXS
+Hh+GygliHi+P8BLvQ9Jh8iDFxVI65thwib5MCUzU3WUTnDSOVzk7O7PC3PLOrLfzKLfCgdC5WDe
hezxnaogbUMF8ajF2M8WSkb8uTFsi02BxDUJM635zNF3s+okUI+0UCdznNtU0zG7jxVUQmXionEL
PT3XA9qVenjOJCHlAkys/NnsiuX7NYKEAehYdpT8qk35f0ZnGtebKi7hV44CADKf8diPmt7x836d
NkFjJ7r2k2dVqSDc8KiDhHJ2pOPCgMYq+yVvsxUplWId6i8+pgZolGOrvXcLtMuRvk19JAri4wvp
YzSRYuWLd5ndQWA7JgAcnL1af4g1/N+L6aXp79fkuXkIc7w7p6kWdJpJsCpbntmob5+ZY//FW31I
CfTGtri+kj7soLBSkOUW29vJXYEam30KZYzUar6Tzvu0BNC/cCFdA/ItP34wndHIu3RmbpvfxITd
6eK0T7e/qZ+KgHF1aL2Wr+E9COc8PcL3rRjVz6WDLTjZ6Wug0dH5OrUjoic3BXESqFHl9jIZ2hy9
YzRQ66cdYD12rIoJf/LfCl7WyG4qM6jL1BoCs1xUx+Xeqrg42/SDy6BvVwu0otIlpW558mykWH8M
M4gWYaq9yN6LeCvgBhDOgnu/kjKxSqrsmP/KcF3rM66+bcTtg6ubppJAgqeLLWxtSVcwit1dOQjU
fpqLNSpcszK1BuiMZ5JcB6HzZwlITK+PcM0fB4FIqAeyBm7IXBkJpuq7hYPz35DZEDQUdDAmhC+V
Y2Oei71YP2dhjRnnni9D1XjFQrxs0XfMKiMbbN1W8hd8b3sI0Pr3fHuTqRFn6CGdjd4HZC9zRV/E
U1DOTT7ia6lsxnAx/LNCatuwkvCqPDTZlNK6gXLH3oi/SA6mvQB2AEn0NkGKU1b3xT6Ny9D/SaiS
WMTXyLuEyIg9QUn7q4cDsIB71pbvzGPS4X2uU4z1WQER6owtFFxwc687GdjpWNfLeebIj1MUE4zk
R/oPol2UnYUEq9dCXV4MS/jpdB0BLKrVPNeMV0KzJtFHWp2I7/V2GQ+wYKfkV5s+Y0Ra8rDOLAQK
eAwtImmvX5xiU5+clRt3XSuzSO/HRgiM9Eay/ffe4GDdgzn+7OzculZp1VMe3TDrPRJu3zHHIT/q
IImAnge4T1wwzHnAuH20UjKejiG4jvng1ocRdmtgudD7p0BbIx4rtjDKotf/4e5qvD+LWZCTvoZr
w4tterizd5kOzCw3ra7EfBJCyenMJnfKi6+yW7aQ0E2uo6nN/uc9EBjIGW3xUUhh+ke2b28TDVEa
clGNs812d7wX3Ii6eyvydQuMD8AdDwAeEZBoFTDoFfQ07d5eJVDZ5UW7KJqn4Yl70Pg0/cqf7Is/
SWPGCr8IOLjURUwnhz8PTVtolIU0evmB2pMXFvHhJtlt6LliZIuoytXYCS08EdtphAjtW92ucjAs
cIRI+qKJk+baez5+9mDBWU14XXTaBQmSy4Gjt+vbWPG60WBchIXdlipHFhyf+UcrjD1DamnpBAmb
iLlRRgirXxYga0TLEyU0kO2iZdFrdsYeLNVhpoSxH+2OuBYkgOsf1BujX/3MJFgWkCkf8BAE0P0H
GQiTRASD4zt64pHl6797QMPpa8y0xmfCx9xCnW7DZ4UlaqbwgcOxg79faEMxI2ruR8hntty4tibw
+RBHxr+VajS1LvEHA2eSxF5rwMORsGvH4B4fVAbcGfmfIVJKm0TPnKCsLngJIZdlmq9zp7g92bbD
6V5t+jr/C8xxEaKrKm0zXJZ/dyDDYEmbAtRXVW6KTo6APNaX8XFWX4OS/oULu2qxn1xeUJc2aWLt
FBZYypBcwjyl3gDEutUejelP6jLbEuUO2kSGr6Akr+I0Dzvf9LrK9fwXQj1DOXL86j0LYF87Znxo
a1Csyg6Gw9I7/OLUzCAKZl+zqWU2LlCV0ze2cKNHVj8EcKoXmXXAoNfIpqUEKg4cecpKP1ZcZ0tH
IzLYaAQWq/fjmo6rea9ZAI0WWXag6036G0P/o/0VgVovt3rY2L53fPMRLog7t7BEwZGg+aWICAu4
ul0mgpu+ab1Om+wbVC4fnMYAOcXdqmsia56ace8yqOaODw+k8vdRw8/ElsCp+vxiql2oH52Aqo6u
JGV7d1V9Xj2LAxRrvlSyOJ7QmzWXLXOI/tXV1x4r7tWOm29p96qR4VXdD4wfkfWjkI3mZYwjRyJ4
OeMPEw+SC6T4a6vd6YdBrrDdGTtHcGO9/096R39cUh1n4Cc+WR7ylq+NOJZ0mn2ZRpc5AFzJIZN0
BA4awhOsaa4ACCia7tlJOklw/tQ3fA1TaxLV8rIcGMPdn0EcwCRmZMNMgJK1F1TTT9cPlOpKZgOR
CHF3svY2J74pAbhSDYOjoJjGhxSAHCUq1v20blmLgU3KjTUioAzIisXJ+a2WIPAeAMyi3hMKuZYC
5/lG52pYJdqm1X2I8JptewsUP4JCR1Pd6g/4OgnjBMQoamzC0DjDVHEomgeT3ZKXgIQmgWBebszA
3OUVni6BUytLtfAIkVizJ6DQXF9JPAXEDyxiZs8iZsQVSeUBiCcfL45d7Ia0/0GLBSO46yTSVYQ4
W3QAs1F+D6JQ+GK9kpY18/WOFbTANqpv7Fbbs/0xRroTNk3LLsYnqHPWheN18+1qZmpTyRpw+vL/
10QKqyJ7mZfOAzQL1HschqtQjNcx6jW638mnEE9QuLJ74JZgOEM6qmbdmmyU6g1lmkrzy0LWXiLw
KzQGmDepyBeGWZYnyoqpd9at4uYQw/R3mEs5HOZwd+uDyO25aSd3Fm9dhH47R8GLaTRNhWkUwCtJ
wuNBJXa1cF4X/Is3I0wcuzz+Gmn3pdFUtH91PCHd4g+Te6q6jORc54fd8+INIlnW6/OiMoMG3zun
mn8+tqs3+HivGv/1QTdkNWs9NU6Dw5P2AvnpnC2/Ufh7L3sGhXssnzbuMxqyPYFy3qZZ0Rukmjy0
f+eTJJRxRW6Ct7qpvPf3pgpyhVsj182qylvSNUJOc4yrXZwFLX/e4sY21Qgw9jhvS/Ch/Cxb2FBL
nmSo5AR11QmWcOgMVEcVggABQA1vIIa2AsetIwUdeDZ80BMv59HDnKbkKuaBoMOWAzD49/rKUoav
HDHvkHXRhy78iRtmHBSCxgOeNImYy1T8SQgMFfcMgLs/hRs0m8L1HH1oe3FLn3SfsIxvloGuZQg7
OoE4WcurLLF+WKlyFsR7HJfiFvBqAsVnQJlGwxqtcmTGKqAkMh3UwOIbydxu7XKUjokrJDlWn7fr
xUZx367YAD3hpca+ge8x7Kd4MMaWMBFmTCpTYuAazrEWdzJsqbs8cLb9uKUSGrQX1J2fuYMgzBEQ
N5uVab8oinEMQdOe0O+vZqYnUo2ydJpmunsQBuc8xXa+9j1g+Zv9HVnXfr8UDi68Qk6CNJfYJ3Q4
cFPqBFBwFwOwU+J8nOLKVqCGigBZAw8puJA32abgAyP7SdOTgDrNu+drkHXoj5hbund67/Te12IR
LKUheALqunCfKaFxUetcJS7jCmXSv7pjvrtPH4X22toHuNrfvoXkgvCfxHzsFUrp1HezL3OTsPwn
h+/PSM8ZqTRp8TLNXaGZFL5Wtp0XakFpcyCNOOor3N/icow0V1on+Tc4hfBcXD3/c2WvV2YrTHYu
nmwCtMqhqqEP/2d/j4XRZPXH2ZQgQxucVQ6YSOUDadmImntD7Wd6EashSFWQt9kwyXwVjn+ZcxzA
bZGAfdfVkRNCMi91vRzajK9fg+9g47G1gJL8brUXiEkcgF/NFCNBYE51gjJJGBVnhe7IsjnoWKh9
olnvDxHJ2hXbv5UlD/9rj0e8TYI0F4StMqClGvAhWVo9Rt4h1DekKvrFKPejp8gpn3nDngDkVEWf
5Pha1yaW49VczsnWfR/8POuT2doE+MR6nn5fGGzj66dBFWd0NGCBe6pN6vUzh3dMyRTwHO1sq/of
OO4pWPOHHCBDpS8DJ1iFnaMmkANRFIWgsFurJLTJ/ZpUxFjHEk/QwYLJ5bHJxJ5ZohxxuIhhlRvN
DCIFWT9e5JfUuTol8cpW1YZnaNJTKvFY54RZdzHAu63PCm9ETBaXqJOj+X6Fivgs60eq+xRwI79W
0Qx1xxr5ag2/Ayg0QYI6UQNeMqW2+B/GLkPd0hbC5VAKlr7W4/yCoTkR7ckK3kYr3N3+LKFCm+XZ
Cw9iw7bt/IW+//VyNsfo7Ml2bATM6FI9uBTTzdORjKY1gNOCjiA6bgNr0IkG3yq+mkJDrX8FgR2/
SUUcVxx04pYC8TdsNSZwl5DPTsYLvE9lDUShm6vvMtCe2orzegoVWIb9hIcxM6OZPTdyZIhvz+56
FZ0QE7YhmZTgaUbJiyBooorp6Te5gx7ve2GTtODn+prOJc+u3EW11c4DUtyRma+H0LLtyvpYTzQ5
XVwWFLoKw6vYylMfOW4cIZND4ePBaTgVOmro96Ef5QnWjb5ucfw//pR376z/gzufmi4Ht67pk9+e
qIy9enct1nxHw0Tg4toHFqDCYbvtqWAVEanSEGZyKXVrOtjvtQ+eBQOdXIqJN55LRkomzmtcSp3l
9kPmAarGngJJpq7m4PEf+vO64vKWhobu37YN71vObtnA3R70tmBwWu7JGR5V9iI2pWaxqyNUk4Wc
ewIH+Z7y27jZ04bScFxnJFVGXCeP4v1w84gsnDhW587B8O+y6oK4mNNujV6fK5p2Zrd/Hdxma41n
6DrbWIbeg0qNstNZTqYjHLWOb/+LSfMTdrDFtPNZKndegHsRUX7oDvg7jd4edQ+KpcKU4IumEC/2
8Jt1meTfAn5cB0HYVRecjCjE1/mvRbzWMaAN0zmQJzztbjfFoj3IG69282zbMJVH0szoDo+zxDHu
uSHo2GGn3p2QjLzdhB4n7t0PcDdBluAzCdx9Z6CVaSFCQjPnmY2V7z3n+l/MZtWn4AkEppzAemDD
cC4Nj7yK3jxSftC+yPjXN8x6zzGcQoopW8Hf7fu1xjnDqxPCC5WRJ2Uer6cmf9NKOkO0pk/EQDB5
/z3YRJueMfGVnB7fuLAOmZ3CYaHcdsfzJDA4t/0z/wdp1WTOaftKsYntIClP1464VGo8VHzLIHfI
6+btuuSIw665tXdgCaoG90Illz9Hc9/3c/8J3FOC8eHoK8n56MjUbNcKX+fm/omzrnmFSgL6KOPr
w9NeVHyKf9SqA4lWdqB55iziUfr+p/0Mg4th2ctzjasbeWki/4BbkAQsljCEY0sr305vWhH0oy5E
NFbgEfeqVHwIrX41JSHBqYZJ3eoJ6VCu/+tgpVAGuU4zH1GDH0WAwcvCVz14eukRNGcW4K7dD/1J
TRlfPmxffYVgfOW5M54k2Gs3dcVpjD0r/Uc9G5OT6IurG9zCNMPEgwTLnzJ+fZBD4aC2ZgX5gTh1
8wxqqHFDpHxm3CRqc1nWOReAFw/YJ8LEVLozctZMQtaVicuniLzGgonTIHJHd9nP/Mi3ndImH1Il
s+fvhDuVtuGQa8QKPbHzEZVTnBLpr6bRwL4bHeRe3yYr1pVNu+6/o7JM2yXuYGPGltI+b45NJAl4
KGKwxaYf2s2hm8FpnT4ZXXGReDQ62m+ncXfZTIxiS8JzNB6yd+1JmHC4dgpkYOpVY3AXepwQXqow
T5HnWs0xn//fHFKuhssHvU4ecLqPuxGDk6DztPoa8KCn9Hu1BT8WbULUi89GXGJU5+Ka+amlPMj1
nqWFIGskfnCM+8NfA+X7d3BgImmiUNFIsz7NhKVekBYCCOZXYm1Df4Ctg1o2gw9KFqx+BMuHWQXu
fUzRrpbJOR8HRBVk25vbdSmziPFe21NYk6AA8jKHV6C/Ha7CNGmMuniX+7P/yPontx5kH+IzIUSU
ieHztitjC5/YHVftEH/cW+P/rCcl4kVzhtxzH1Z6hpXAmzgPDvl3tpteSsqoQhSfuqSNK3QxCPQc
yQBbvqwityzmSODn4Ar+wD36TagAYpl1cZxjCtmXjQG5USt2kj1vWEJIVg+aPRnYwiRZAVYoigWE
VStnorNGzx1o9LGYeWATFiRW5PraZNbVxXWmNJblS1oUAZE3gZXLkxsw9wdyHMqFDmWmDEy6nczK
CYXE2MxkVcSXzLnDAqjPqnGgcT+VU0J/pwMWZij/dcmFBVM/nZC+k9y+SdZqKq6qK8E2cx8rWDdr
mOP5LtDD+BT9A2rFBmKTIgS3B6HAyfEqXvRWSLPVHtNanXWBwb6gSnECJ/sbsY8r3Owh8c2XxWa4
hGfzOE1Pz+eDDB7oYZQ66c4JbWhVQgk65aGGCxffLgQqwK7YyOgG1ovLlTMoa2Vtembf0fbmyguX
kMN+yobAB7uN8J+xU6OBvdhjmGPe9NJBpbaacClmFI1LfFgPi9crvqWgP+NEaQFbgWb+C63krLEJ
2o8NpN3wYHHTPy3s17YKYR/14dZakgMpGFUWGCCSIysGZjrx79AMTRS5BoUI8SIT6k/ucozJ4aVA
Jqqq92QpzhK09EjSS1OjWuMFgIcHW8vJZfpPdRu/+SgsZ9oRcWzAKaDStEeBBBI460OPEVMIdrzT
0OoKuW76Y+4koFDmDSiThiQ64yihrTkiSQGf0YPZFWxeOwH5Vxtn843BseMaqE7ZUqYIudPCy1dT
fWNqiArCf03gqkAYZNeNu1Q1cKQ0q/ofDPAxRCTXbPUBTVqrUPEuw5Rdqj2aq0NXzk4394BllnrX
nEh5F3ATnyHe2DWwUHuBLiuRUDvGq16YRnFHVRN/Y53WlEaD7Oz0bjA3iTK8bEbXTO+Cf/pc6EKo
3e80eHt7mAkMIWAdrQdA3kww7ZPsVXamahgfOqDD9bVeHgnLG84fGUy3gMwiEkHrYSj54qJzlojt
voaoP6nV0U/Auo/iVGqaDdvMi5mhxVhpyS+YjEQxRZ+BpAap7BYYxF0ak8HrjiPALlaT5ru7Drrk
+1W0S4e/z5qD4n1/cDCmjL8xzvgIJlVOw6ukZGwvBc9JWETIkqb0wdTHG94iWdmkuL9lgUnkxQN/
eLl/554bSkt0HuBvoFB8+so6AbQabY7RZbBXqljl9ckk87RHawocl9DvrxIqa8PWOagt32+yLWRP
cdzxKF97KJAli/eQPrT03B4F2CjIW6tWAsRe2I+Z2G7pee6xYIg+ryxy9RiADtp0S7yvQme2AR9a
eiTExFqNxPMkcvYfRtNy3g9Laveb2OT6/JWgK1ys5bmoiVMyvAVQ28Z4pYEXvO+mPjb5yKnFuxMq
h3eOtpIh4GVS6QiEVwgAiX31/AHQBX13BSAc5ub4jqQQWWe+tINNMJ2yyGGXZuFerbkog+odZwmh
XuGrHAYGsEt0MXB7CIKwfC8b8RRwLRwL0VWXylIVNNuRuJAtwRAsr7UMsXmZbx/fUK6f6Leh7sfK
HlM8VEiM5yyFmkqAiraBI2McQd+hrXJjD1acwU+XLUAJePmzIAJ1pugCyJgPdHP820yC82ajaBpv
a9FwdY8lcRLXmNKobR4P2gg5ggheVP0PTHMr4sWhv5f/m38FCz/mFbk0noZw4JZe4U6bo7CGWaf3
heXjoCqrdDHu7j4b0f9FfUaztyf4lsp5coM+9qyQw94ojOlE/3PV+AlILb+OhEbAQfeErAJZhtbg
FZpOK3RxujnRAI8Xyo2erZp/AM7yIpTtyf/ObcSnzkyrTntN+iC3T+HZdBsCXSsDCNTFiUnwCsg/
H3SleejbEdSFVa9j0ocpmLPUS8tJH8SBAJCr2eeYcB7tuMu1oO6zoo3so5W90YjPknE0OclOQgNg
Aru/+qw6FHqSMkKLoEt/ImPrgE/emcW2xSHiaoIK3U8YHC0/ADFDix2KoA0pYOdcxjn2kMSW4YSE
lJ5imgOMagJVWNvjrtG2+J/IzLYisUChvKAV2EFl4ocQYkIfEtgR9t/94YNqFbWHUpBhyqQTzy4q
5gXsZEp8I8bjalMEgwmfueaIl5JxtNWZPPOuBnMuOw4nJScDomskErvqz66OLFe5HfKyGDg9WpOe
7CG6qpqIGLtqprP4NJb2mxv5OA+G/pDD+SnFd5wX1LPvWMMQjhpKkEbzSuUMOdbzuvPsudbF/p2p
+DGeW8VjoxFfk8uZ9Yq8kJFMW/qTI+T5CTohkRbhznzhFZorzyXRs0FRvcq7kL6zbPESeAbZkw2M
V90bMb6cDAsH3EzcILSBc3+cQRUReGZQ6hXReB67SHuLLr5Txv1IbvqONI+DF8UVKdvOhD7FwalX
Gg/oqOrYZTfc8mB5eRy01QUmvJuNFbdxLShQ+oJtzJj02Q9Hh1JYnUULTsTKJvMvaGKkwDMWUhkX
UhpIFOgSiZ40WX5zIRHqNvUyPWSr3QiA+F83krChYEznLRPFVPd41K5Q4+VXMXEzI54fKfGIgZjO
GKBj7h/TBUGNA4/U7dnA0wIN/V3EjdbQliSOiN6BpMo0+OTBmsJKI9FXrjDOxxWOC1RGZMfW2atB
elC+QQHwjLiC8yTbH13BF7i2DfIukyjoxBoZiDcS7oWGkBz+zaguVYIg0AlsvGLuicmze33z4HTq
03gdqGlPsrq4/aAwRkeohrbbhKUA8H7BI+hiyx0IDtDlc0SXI1lpD1b5nEjjqZW03fUIoYtFJCxp
Bn6D5CuCjnL4VdLkKqHOTJT3VsHQXqLJ9Eb7fV3rj+xIqoHzKf05RtujG34LfN3Xt5jwaleycoI8
5FIrkaZSGnOZ/4qF5/21m4MPjXGXsVrQkzVZVZL7sdlunI4IYS/EQCei+IpzsNkpxVWi+P5AwOJe
zpkBKcPSKsi82vehIQ1DeRl6nxPwRKxgiaG35FXncH2uMAVKaE0b2tZAPg1BnM5jNZ5NlzSnt4p1
1NayS1mNWLjrfngNcUN5PWu68tSERfzYVyshj/daHyAwLjA9X1bwPU5+Nw8fQCaWE2w1eTr7VcqZ
L1uu8nGXi9zZXCZ8G+TqM7ZJnB6294HTWJcUK2QkEUbKYOQ+W70kRinlRKsIkuIc/IrAN0blZ9Ar
WHJz2nD4G6v5wBdeG8ctgg7wTiRFwUf6eYjoGymBHbt+sh5UnftxuG1vK/R3d7JbOaUc5Vkc3kzn
4NiS49XabHdEuhEx389g1GBajfGOct2rBUrfaDkO2uhnaA0B9CBLtxWf84TznwkK3JKLqOKN8cc3
S86Xv2qZpbWhf+39rbCTKIh4MPHyUdIunpDxIDZQd8rx7ix5Y3i1mQSPSwmEaFS3IdT06RVlTlGE
OhBy1feUs6EWJoqLQKmbBGHYJifo/qHDcWbA8ulUghnGy/xgp15MXdFVKH39OzZp33JcXtyyMCpv
5YI8K4yLIt3nDr8giAH3g+sgd9yWGDTtUjw/FOVygoPWni1uSELmktl6xgf+8buypEiIS3RkwM2k
aux5oLLnBuYYf9dEpm5920PDTUuhxYE5fg77In8kyNzpA6BARer9k7/ynyh0xgE1s1+RffYxFSNw
24rBmqS37JxueVHaNTyCkPnfGqNmKA7nV/5pjNqzeZDHCnsBzsp9cQEsadiG9hOGwFopfwlA141j
ixERUO1rEHqlFIoTIaYmJTszi0d6h4FTg6qrVmwW9pzjgZv3YACrHavU6o18LeMSTEpP3G2WoOWm
Idn1Lu7hCM8XgzIDwU5FjzEmsys2PXMAioEK0ce0HAr4O5CwWf+hIc+KD8b12ofMijn/PW+JhSr5
rhi/OlommJF876YAn/LAJtOszMbYy9J77yliRGJq8ZHWKKctLoc6LuM7X1KmbIsp6i/aMDmLl8Fp
AT1lGIWly5Ldubz9OJCpBTp7AJai3FUE4ghZWzQWJ6lC4UERF7tmKMV4KoZzD407x98d2P6GeqAr
67gxExU3eMzwIL3qtTNAI5tvEv2vB3TCx6dQCpYxYuSCIumNdwy/YZ2XVeNIenQx0/81xIwnRhZN
R9f6+MCfj8/syhApfmvzsNO/fkChedK1qHRThI+x5Kwffs4AF7xmcWfb76C/PquhOauTo1e6vHgs
Hxz5dgy0QjWq3U6tz+eV9AVe2Xccs2Ug9Mni9nlukF/zNQ8m7lHIeyACGI86ytRRdXxciiJ3HIqh
g1TKyFo/pLu+LOL5srDSynP9uTyxbfH5J4+89LA9RIuusIl2pVpqfcYgol/XJsuEnM9bkLlp5Bwg
idlx8Ziui3ZGxgFh0eNgmej7cVHq0ALtlFUmZ5NxYJ8AoGz3LRWyuxwNCFgV96oRFUY35hJwlkEh
S7t1LAUs+Z2fDCqZmmAPO9mwebbWPDRIipXrgumyit//bHkxgUHcymLbhGU4d+BuUKdTvM3aamjp
y3yJRpH2aOpwtWXqllkRdEnPbDa8jj2oG3qaAVMPjnCfsgxKwLwhicmrdzT9nvsDxlMVD89VqOs9
SSGvxhW4R0AKli8jaoWbgTl4SHf27H/y+D2yVC+rdK8TdHUNQrO38DbhSjNbpAfjGSN73bMw92jA
KT0/aom79AAjTRBtOyCyk/LsxkTR0WpHr+1WVpvJCfkz8rwVGh+Y//fwLSay6SDSHTPgW+1dqfFy
kCLYGidqs3EpMIfJIBKIDriMVHJ4OMj3ODjoQkiFyREexPiK+oNmCqMf+/t49NpJGXLkwR2YJ/5b
4hB1FSfVDnkPJR14Df58D3tRXqDw2W3y8AyqOgduyNpXIkeb1RPEVNaPUybN1zhrWsir9JrrmlFd
khAltXHchUX/IzXbl2hAeDrLR3+TKQAVi99U6Cst5ek5A74VwouOZ3fJL/wwXmMsaahm00GFsj1C
09+p3PL93XiHCeAebqH/L3nsjmt/HG0ae/Hx+kxqcEAB5dJVpHqqSgAd+YwdyWZth5Cb3O51qrvR
dijITRrini2uzgFanZ5MXY8EzbL5XTDNn0+x1eRBQNpxBRjggyL2ygnXi6m4ImBCK3R50d0sHV/3
YfukulHEULxeQOTUANrZQL3TwtPZSLm1EJ0VYZfPolJwbFsF6UVec7Y6lC7yHQkbbb/tQJ8SwoQJ
DIZ0Ul8IkCDa+Af5SgstawBCAwsjCv3BgcEaRWik9DCOkkbNPAGhwiMEAO6lP7WSImd7i8617brt
oyxP3BsJXontY+I4HgF3T6aAkziOaQi7f32JN+MyoDrkX7c5x+d4Y0iKq8zvgCF5Ot2Yf3WmUTJo
Oddrt5700pkSB9NrbWR2c3D2ByCwtnKDASb/cVAnfe+X5p0i5cmgwI68kGzGsc81Uzrl3lEk80v4
3DetfQd//J/316X/EI7PSvNNo+iF4cLcu7zJ6qhwbe1i/NkCmnBSmMoGErI9mTycQNqdiW6dW02g
7VL5NklCEPSRBupjP6xYo+LuGCOtYhF4lcogSY1Vc98rfm262DF6RayLZRcdMaopE7JA0Bd9MfgG
4MUShBtJWUw0yODCD3NhZeXfFPJuXc+QELyLzq3diAqPpwp/kDFARMALBQ5fZbZp5YnKLmSXqtOK
Gp5r00yEDR2wHeXRP2AVPBz3klW7L+vhiwPQHBmSXNwOkhi+d99CW9rjx013iYYCUBv5D8V171rS
uXaxs3aB3gXujFQ/lFtZWY2jyZ9Qr98dPpre8Sbwnk5lOqm1vggmpGIJiPcEd6BqydFMItwoX6dE
6giNCAEXSTgbMkNFcSCPG6C4Blue1T/ON8IlvaXMDEwtO64kyqQhBUbCeRDitQ/aFdsE449PS7pF
yEpcAc0PPJJQGy2Fp1vTR5R9YX3xVRUBB7QHXOzmxGThmqE5UZP/oHnrzwENHV0+vqYs1uJ8CQ0B
mKqkBthk5HpsSMpL3RA1nQSR/unfhd/T6dzIv9QbUxXULVksMjWPC6uGx4241YI1iv3Jb1oO+raq
K/jYW3feLEk2963u5rL1eAdXSvPh4dtBdRUMwZF9gfv4OQ2VG/0Qi10nI0pFakB8B8a6JPSUl+c/
vrcY///BA848iTPCVhukYSOElSl9sSAshBmC9RsM5pj24XIQtDB/OaANnu5QUHg5VAgI/XEs7ano
NtLdkjyXxYbRE05A8zKGKXNCYmjrT7w=
`pragma protect end_protected
