`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Jo0GTP48lurGV9QI1c62RTUP1YVEamMz1VZFzIOsgfj+B/Me/Uz/+TNhvOgX00Boh3rVDWY3miWC
6dvD9WUK3Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LQaetkHlTEQ/O2QuW4ImDf/K0WBzrX60Y2eOh0Fzlit7V6+gYpu/pdjpcV2iUJ0OSkPSJI+Mhtnw
My00nmvcw7hr27JQMftgpSq2KJTPiuvMTKQgaTjH7G11dDQzZg5OIfVuhiEdrvLjBL6ODFpLjnot
+wtza061w0h0SULGF8g=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
e7yz9u7SkKHpUf45ToebPKpSB+7SYjKyIPDWMVo4RpE1fApRY5i+m6AdkyczFN3egPL9yuxMUBQi
B3fcWe1KL481lABpqgSqODHUHO2V3VOpcYtVbs+ITdbbKzYLqgggxX2OFaFxfaKpm8KQDKkYwb5s
hDH0bmxkegiSbK8/6cCO7THsM2QEi5MCtiINLnSFKZxzW2n5D4XuM/reG5kcwrmcvNmgwL09iDms
zsLNFk+KlTwGLQ+sjNp4XMp3wRVy8au+yG/ZaAjv1SaonTr0s0Ktoq7kpKzzK8Vdx3gxl98oC7lG
qI6lKENHTJsj2Et1sJqARwUVTfXhIwUnx7z+eQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YUgiCLqe/j/NhPlORdPixdVwbLBtEL3BY6gCgf7tGi15P5FTCSoEIKV1fMOt5n55kUiULz6ixyOx
w6KSNkCTxNK1tRyjWlYPNwh+30X1DX2lqxQedujI8dEfW4TThaFzjbr5VzZ5Xx3QklpDtemVWlfc
v+85sRR7dpK2+yz7JHTpwsBUmUIz/yQuKTPH3TXkcTEtK3SDtuMd9W57I7EJRQs/QWb0HRC1gqri
b73Bznz/ITOHvk6hyVhz2IcLVxpPIWw2SPni76CtRBGxpvEkYBsB4Tb29iojsozDmdeCBCdMwy/R
z6g42MtTw4HdwvXecIHU1Ps+g//YLogOmAG9jA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
m7rYtXUavsevrUPbAA9ErlXCOGGk4fAoeRrucNOvvuTkTuigciZtMDGFuNCCP84AUenq7yf+knfr
YxGJdpaWbSksXpHqc2OaU9JxiGbOYXsVLB6aaIcsBViJ1Iu9Y3dsxqVRuEf/+KOaUoj9MgYpzlBd
dGJCSN02BKWDuiELCvkTzxH0HkaQw6L4Fs4eaqtvZO6JC37ps+GYsLvCsUVOUrxP3ZXffR/5rO+/
r+Y7T74S//4yP9CGXNTnVBNea7FKmyEzggzbDLVXfwg7DC9jqBdVLhJdArtJhH0AWfbyCLDAfF69
TIFn/nOkcwqHGmFmfhdLuMOHq1GabkUC03gqCw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WkzTVLle3kbJDg7jpvQ16rMwFjgKsN6s5VraGMgY5PuWLmuM4CseW8hGJcsf4WjZloefR1XKRkv+
EV0MnXlsj7dM99Z1mYpSYEt+FSSlVw8ZrTFDfAXM2tVaQ6tHWq2thbcjDszMiCZNwxeaVwffojNF
dPRWtPW7gJ6hRMZJ1oE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nB0LvvHetoBgxBsMSEPN44HAKokSVtsq+whVeE4wsASFbqJ8K82xM3hbmxu6ZDYkwRj1/AOA3HVk
G4ilfKGLy/G7TDbQDfRO+5Y01cbhrcP/GMxbBzv8olyMaD/JTd0uTncjO8AIV8tUE18Kj9ZhfRCb
zatytXSeRs9JZ1gbnMMyuS9DWHly6IquSzk4ICOoWWjyjXwHRFPGPkYHKeAKIXuBgNn5YIUb73Bg
ZfSxBEDnDG4lR9r5BsXVWXPmkRPzzmalgCEOM4dNamRFXJG6Z063apEzsaFADjlPswBxcO39daPt
PO0nWMUFnDtLtq5NhL5JcY8vaGgEnfVUj0929g==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kx2/4FUG+WgpOeMb3Rbb/cih1lc163wBQ4vKkckklmR615Brrk0uvh47GWx5YPIQIJ1dUYGfGof0
suWssmlsLprBF4iyZ0oJN+doxvhmSoNuyqNtF4sOBh2mA2fEVAiuuRzdRQMw/lsxuNxU5tTeu4Hq
m6fseqlUS4i/DqAjB6NT+vlMZPYsrIaV5xH4A+ZthsSp/Yv1VhT2z1Yf0I1zXIDSJLePBat4WiXu
ztJa66W8SRYkuIFjEUecZElA0JE2MfS3tIGvepvw+Jw2NqcpRNOyHazWtDF1qGPoplQ2+iAwhvFE
swC4IvCafgzOO12FbZwI5Wi1IC0+7hrnR+7e/A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
8GvLC41uBcFwr5Ki5OvQAwh2MwnGKfuE0FkJhaohC6KDT4SH9pKcwnvFqbHTm7H+kxpfjlg3NYlo
R8dPW4XArskiR6Di2uUoB/KHQZgA9Q2mfXzTU8Fbqj0lQxpHN6gq6zFU6JHgsXkY5xw9NuM8/MSf
6ADEPnXTx/pT4gaRbv58Or8Q3mqS1S68vZedqXVbikKdIta94c4Eg6J4Pf0rwVh2p/VpONb+vi95
xIIxUGW0no7jVOWO7k1PUT42pwqJulTpqVAWl8RpLUs8/7LhQag476lWpcOsCf7Q0bsXVbUT8htU
LNLHcGfqNOwRPvz06K5luDpLD5KAXEP0ZUFVU/YsCK8rE69/I1Zg13WW8jVZC5tyxzhihgcNf/rm
EurloBPSbpJ72G1HHwjCI099dbSDlDZbUJ63mHrZKJ/CBKnqODZR7QgfHqld97g8J02rGoGzof/m
ArCXlxajul8n3jXdTjh6+dwB5kwTzUc+ScSmCF4sYpDxtsdezqq/ELRxq1fG45LIOE96Y99w+hQO
IyrD2FwK7p19AW0GTPA+gDfGYOmvGptZwnWKkZd4ef3T6xWm31Hy7DY+zUnQsJ6Q4gCAxtQZ9kpv
NAIhZss2Fu/T94BBJfZfs7W4ckJBFqPYPfRcd2lkLX6uu+MRsF8VrSAqzLEO5YsD5KKxdF6Jxzb9
WnpygGh/wVcqrnXmTi4GbHqYXxu1m9TM0FuY4PXpczDygChfe2fJ5hHLG36YkbhCeOp8eyF6UnqT
mRcm/KV4QRIEufDxsqc2yLIrCSA6Hvs0iaLmin0ROxvA8xUsZcY+c6Y4jafYysvClb0qw2dlKIh2
Q2lpZlPapIPxgpzvPIFqsgbF1dsuSpBOtB6HAH7kRyZyODZ4ewR/ii6x+Smjpu/Jcl0hHSqi+zEW
rBgNw7NIap441LLZ8nURVPr6ak/rF7m4IQfRsDqSZDncO/t+bN4leqY8Ai6N5DaxmsAK4lhrqFV8
lwrKvSajRqEvZKRxc2LFfNFz7q7rApvjKl1MuIaewJJa0xAysZA7/ZX4TrTljtEINQUITF1m2MOB
q/XMHGyCBTsGb01r7Po87jCOswYcZ1TZLqIQnifvrVd76ez5VW9wpLuB1vgiFflZ0TdfzV+UduMr
8woCayw+fL1GQgnwdbPR/BANf+MKO62Q6VP4p+amOah9dj0sIs49+JkSXzCuOQ63uRsHL+On3094
9AE+jk1G2XhJAWg+CgI11rMGIrW/lSvNFKgWbQ8VdUao9QGOHTs09gTD5e3YUaOKiKzpdiMeovCX
yXeF/+au0j/D2vF6aM6tYus9QNT3DtLMI97YobUmoM7CfghHmlYG/MwkAFjBcxeRqP0IjCpI5Xid
IPySwtcbEHlzWbJrhPu/kM5NaAovJuGDALoD90alWxr67me4GtBEgmWl98GVxyeUyXCiy68jw3Wz
XlH67Mv/WIN0EvatrOsEDb/E0He53dAYqss4jIjzBpQrMyt9PYTCvB42PGcB0j2DsVy79CEoDGQ0
6Dr4bryRE+EerbYDBETSxL/e372+31cpaWhKHO0InXbnTnCQ/iSC1Ytt/yBi+xBhSHAbWhPJSAzu
zOmDCY2SkuV8eftgnmWX5STR+Ou0lV+J+TXLXFi4j9ZlrW3+ozYZcsnzZ/HL4WZxHkZn0NNx3u19
cCyntgobySqahHW5Mx4n4Y8SNVBBXXGIxVwXamS+nROotW0N4K+eGHsMXL4DbyI6U9dpSnkaiW3a
hSHgjCE2Gd5L7yAZWngHcR32dFalaNIFrafnIYcO6I87hZOtknPF8nPEwIxBl7agnmA0IcafIbs3
duT72F5/L+6ln4SgLo1Zz1hPjfVWWbqmeVpSQ2OPhsiBIpPO37Iqg3FiWdutaWud8UjnM2pZdfDY
ZgSFpWeUjpThqNJyP4BLtdi0m5OxNxq57g1+sYjOKpMZ3nAsx2FBl8kropm7DnXw29cCt3kFZndL
b1+uU/3VmBYEisf4oKUAq0w+QzW23A4Z+EkZ08s4/iC2GqNrdOGs30yChLeSp2wR3pF2excE/Joc
FzUnYJYeBy/xu/jY/QoHxCOQF5gk68DXDanKsqBo6VEL5ItfuJkrwqCJc3pf+KTBUSYuHNesGcj+
VcsLMGC/D+YO3qR0dMy8iLVkr5rF5RnlzI9ZMltM5kmFCQzkHt17wd6i8MiChN/NUTibvBO2Exi8
nja0s5FWrVFnKEr6rYghlCWAFGISowOHtk3lWQDC6uxhYqhPRbDI1VndGeZL5O2jEZYfLLy+pa+1
Qxqw2Cr7pRh5uMQdO3D5HO07/S0R7U6+BlQ5agPawjjuRcSyyLR1xH7SqlmlypWZS2EUkhetT2G9
C/fydtUiHCT+F+t4JsEshiAk8xP6FN7zQjO9kOZJEMkjKAYwce9yU9ReTMa1SwEiujBN3Lcj4Ps4
t+xEM0OCV7oPZfr/rZI3XXjILWdnO8pPjz4/0EXIBn4LiFckq6Iamvw36i1i2p2KbyIsBsKIBfN0
qRR653jUqHpclQBTslV7bw2f2wiFv7irQQ58taLs2D+FI9r8nngCQ9EjzR00SdkTwQ0+X+VsFMob
bn6Pw48Jh/82MSyBQDOXPT8YP34FVrqm/SsmTeXIxyPhWvuisOIE21bSu1u0XD0NlFkceIpohGwS
MVmMdklVWkd3Qf6BgjHR1YkHXR90kNIcolXI1hjcNvXqiTp/0HrwWRlxAY+3s7Uub2Vufig37s7j
+eivbIA6pSRq4ye9mDBnPRvC0+bCEbcrdidHohO2vsuqQml6+5zMxGtiof9UyWFRLNuWdgfPnVSI
fOg1cIeO0ZbXvhoqV/DNdT9/M5ByiJE+7dKbX5y+qIKG55vn3d/pzmUrN/UEZLSnoU3hpXvMA5c5
3X0s52gWdW58VnpP3H/rkHt+xUuD3syn4ue9BzkCqKz56j7i7OR2sURSXFjeWV6vU4RkHnMxU5f/
dpqcyHBH1J0/EnQcLm6reFJ8OMzY7tuXhgghAVq7MMm3T02V9UN5dMGQLiSzKZoNmdqT4I80PkSy
nOF9ctmuRvt+sy4wfs0NcK12aMUbxlCrPhlhCRgv7OatyAzibsrLVP2Rar39mh1qN3TKWfalpdwm
oCjgmEAT7cnQoca1PfEEu6z7VVyfMLXBv6k/sR19Vx8B4QpQQnraRiFNwT65pW9a+pSVA0Qojfyh
vuD82pjtHdP/BbzrheVnMGAU4G5A1qBu3uhHZvUde6A7rVjQ0jN7K0KNU9d+9a7vyzdpw29AThGY
c7d4JSNNBxZ+TvCkaNfR2kExQobRzHyujy5D+Xl3yB6nzm6iA6evufBKWpdBNfyppbeAHp8UsVST
MoTR4nfCQowanWQWcyXGnzoxIeTfx7rU1vR9yOuqovjG3DBVh0NFt+FMnx6cJCn4vXJzRo3M5c9x
r8B9DEDYgltmx2yrAn0TuF9tSw9++/YHl4YdrRYzuhxAdHFnVN5Jkc2iFbPEfJqUu21wqNh2bB5w
p8tzZAlBjLx6iNDRw2ux/29KOAesrRItqJPu9dW5yv5pAxIkJ/1Cv9q9cNCeVaYn8GTCPJSxJF2F
UXLL0/5Uf7T1c6E75a2YhizbeLGsk46nctPl3ozYNQIlIdgOCgcMIqI2i1+reOoWYAB5rvmXxTlJ
myzb1FB5gNZ3bCZraShg+4Rw7JP410+7OrdJG2uV4jmWz4GJub08hj2qwKYlyMvaFSZKydiiimMf
uuZE08fRPmoYwfjiJb8lr7rFDQPQex/6dXDyN3eeoYePiiKgMVvxFIGrmDTc86MuefAYXgv7nM4x
2KSbqTNIcL2WUdHjRTm2oMwROKuqmm3OwNPh+gceORk7uWWR2s3/BBRbwc37pmOQhVyPKpvKXczw
U7xnyAnSHTBjImMvJEQ57r3Xb0MMs3nG8Nny2iCj12ymk5z/RafAOcU5RlhZjJ9PSIYEqltkDebE
i5vXwfMiAYdJlzgRD8WMZ366HsbOsvqw8fxubFQEYwYA4kUXgRPY7w0EEQQji/qG2qzcvvZVLVmB
mn6ZgeRu9OF2XZSBmQ4J4pgT3FXydHKRs1REkDwNJtm5GFlxflI2dAWWMNGN2LR0lB6jwZiPvhZY
huKiMVwUOF7Y5lfqlb504mQub1ebldvGk5u6ysuNHV+1/G35DZNn6AXhFkv4OyOuhsaX7jDMKCdC
/MDbArJzwoXh7tTkQYmkrtJX3DOM5NeSlmRRSKchsWjKu/a1cFU621tlUiyFlNeN7OBC3DbNMwxk
uI7ecdksBOJSOPHR+yJnwrKIqzYfCCECltSFB+C+qqUWqJCloHHuQ6OxBILqP2OfaPTiceaPF06N
IGNu2qVliTPN4CBNWGK+E1Ak9zMOrEJsHnKwts+xgndwNCspxhiTMXa/djvtbush+HR5uhdKfYv2
I3XcDBo6m+847c4LsNxLhXdE7IvQULst4Vr76Te3JmEaXyM+SS5F+vSK/R6QvSUEpNAsj7sj6f9c
GOucjXO2hKS/JhID1vhcVJihdR8LlEWVW++n586aQ3RYt3UgRRaeKrpHPXopOGn/gj2jb9Tt50QX
pH/2a5dUD8wMudI5kMhQBeBDAHYteeC4mnS3BWTnZraLWK2RrQGFCm+H3/jLFO/jBnXWjoTl81Z9
+/K/kw+EoqzFdwdIu6c917TlZZlf2rc3tt6FvERBNNoRtYkmw1ugcZ+aBO962e76hU2W+PXEvZvC
Bo+RtIz0ujPROMu/ewrisIOy54EKx0ctkAImrGZZcvjR8TzqRTRs/voH4QONOjTgFrxgS90lRcIl
gZQZyebsZE+Ts6/HIHXfVgsOVSYthZRJEcbYqs6CSD1QUQ0/c5IyjRqw7vNF/WgA6bhWeS1g0jmy
j5suceE29BBVuv2LhkfFwlYWvIfEKQIi4d+qMxv6UVHm1eS+qc94PGASRcXCq00HPfwS2FV70iTB
ye5yTq1FhhT0QGYxjyHoD8MI3OQO48dnMvwn+EUboJxnosQBzb95fhG2bMeFMqr/Qn9qTF9Yf63A
xFA3GvCSFK5biLjvR3tTAq0TlZA0TCwMJntVR/LW513mAtVK63IrqzJJWOctjLd54NpfeYkLnhLX
5im17VNUwDQTpsmt3CrC95YmEaZc5i/aHShDpg1XJGWBENM5RLVn6PLhVFJP8T5M7vxRigU7XwZa
BDTVZU8BQSi015yfgYcGEhkYB7w+wucHJST6l5hp3TjAMunQ9D7G5WUMvkZMYE99Hkk4WM1dTLDb
SJPAyvqlkUjyA8fkgyJ3YNasKuNZGVxK6+iY4SegfNh60i/j31kQirOjNDVMwh25TLqx7ob+6qxd
jTwcl69f0w9MfOgyzysQr95qIfIwfCqpOyRrOrDDuqq6fJornm97xphvkCeD6wWWyoTI75JXZByp
e/JmAHOcs59NIAkasopeulH/15xmbqQWeYIeT9htvygLYV5YVjJAE4FHscxtyBbY38CZb21POFPR
0iWbVAe3nHzq875gowqLLWBVhyLquy4/2SH+UpFuyitmV35ssVtkJ81RGUl1OkeEYE00vJ9I/IJR
BfWhXYDcsXDUOSAmSQ5PD9hx/wqwHS85dUd0Pn8iqrj4UZqOh/k9l1ZwyN4UGAgEqgu6c6np5loi
yk89s1sEXao8g7ZK4mZ0U8g9tPJ/dsFOPF0jL+MJEN5sSUVA7PdNvOz+CVkzliEzDdU4xl/jJOvA
ilLDIBmnV9p4QuIHJRhB1vPmd5JUxp4t/IA0M+44HqSCHu0JPR6+FxXqaZPHFLn4a/J1QLFAruoc
5ckc/JNkNPjKzT8WKHknQJqYoDgbJaRBZNwQ/00CWjIlIiAyCaHlwF3ABVNPjGUqnO0llLeoW+P4
eHnW4GHM/Xhx4I7EOOkDr9Sks7CleRuK4Wbt2fxZjEK6RbIHcGNKwcLtOEXDmIf23UFbyNFhkVvD
qX4BsXUnc3OitJglZgc4Nps7id+wTxQ3TxRvASOvntoL5Hg8wJY8CW+lcAXtLkI4iBY0B3cc5h36
nCMPdFlsfYWX6IuBYku0Csxs9RQ6PFp3zIimPHne8HCap3IQUNuI/lWJvNKEeX7lSFdlVCl/SBlI
wy38+LvYgtIDXX3PvqGcvVdVsAS66USLFhOV+fkb9FE5C+n9HZuio8Futrv8RCXPSLA12A8oeO2Q
DH/O9kTlFKZiUVEqgKvCElIdDb/SAGsK3auH4E8BnNhFV4ocTevvwlQFN4hNMScFtokKWcT5oPu+
aZoFTsqXu2gUeVwER9XnjiEPsEoiyFnhdMIQb3gmdVAvJps1zY3IFzhfZ4JY0BwsZ4ZPdOLvM7bn
O8uWd+7HCiSCGUTSvo0kmE9gSFjVoxLWxfLyBOUaU+hKyf44ONHnqfS8jU8RC2WCL83Qhml5RsOO
g2Um/rFuaVYcvcKQEqEFKyBfxmYwXI7XzIjcMu6jaO+0c56/savcCSS1qiERQwebcSayNhTNSNHT
hDzGQd0Wf1IzoUT41LEf80LTpv8pcz6WMXO667UKOlBZT8NuTx3cX2tJCbMxf7drMiOSsf2r87D7
b1sG7tS5MIV/73uTeAfcdZ65R2tJ18Ai/GCyrqy5h/AxqA8Z3vDcBJRqvGbv1O6qtSDtSZuOcmXL
4Vsti8pIyDBk8PNB2NXvwvssHaGxxGOyw1W3Ozu5wUG7BCjlXxfPcmRlxotW/KaRX5l9fDQSm5Zk
3ilk3HKaogOPMuumaWoDifkTH7tD4FNn3xrI0xfn1yYsBedA6k+tZnEYDCPwzjf2GfEHZ9MsfmBa
RqbltYADlrvR6MovBeLCc2UC5/4K8itDVAxHWZ6y/cBuW7nDb0hNyizzy1y/LmPqC96bD4u+HVuW
CGWgRipWgqx9SYTSQ8yS1HzYapHfQK/1W88RXUJqTIBjfBGpV1zCjNp0yFbz5Benr7rpZIosnvtF
YJkj0HJ+7VXwIeyKVYfTvveFdJt5LGoVK4vfz3UYrx30S5nKrLSUko2dMw7OkQAYyVhGcPJD9+8l
LR9vE5KoAW75fktbQ89TnKjnPlc4lWs6P4YztOQ5lDe48itUObfI9aU+pFJqPXbLfInMdHR6J0Lb
LdRDlat/KOJGBS0FMvDDPz8QDoOp7onznMTdJrCUwYcRXYhG+OClaWbsjYbegaUOc1Z72BHloUxM
2WOHsm9shtBEXCCqXM4NMJXrYWRsbL8pouUD1DiC7/JQv0uyisQhFlE7QfWw/sS+T+XZZNQV3iTQ
a5Lk0EFVbdL+ONpwF8CoNcBNiW9yN4GiP4zb4VNqMtKpQpQbJWjn5P5TSm/QL8tY4meU/W/RaP+g
pW+Az0Ac9oVijnw6Zrdy+jfrfjBRtrIJL4E122Xf32oWFvwgvSvwZTt4PhLrKo1oYW8jTOE83YyJ
8VyFLr4pmuFQj2Wpf5SmWm6XZvlsZCgAqvovwd7CKZHY0GqVtscB0W/Bp/GQRde/qwivBdluHwv/
ykTdapfx7soscw+xiHAea7hOBA1v1+Fh1HkXgyNUzDteYPG/fia77VrXjkd9vanztH7tRaOxFfcP
L4E7XZp6UCaBRRliIoPLFO+ng2P2YCvCtxBHLKcJaP83b4Pp1HG6h9sDhbEPw3lclbTLRFll04O0
m3Ov7eGS4En5T8e5nPjxtZ1vp5RrkQ1cefqJOJo7KxehibhApURbnMl6mtntHzCWlMgT6HNZYPZJ
UE7z0KfG5p9sY0KeMbL3VFCRkYTxObYUJ9CVQAiN8m9qwP6xIl5hVzUe4/8Hv0d4ZQXBX2OWacf6
PEKsfdb5Cn1p2BC7G9ctTDo3lEACpiXMUa/G/AFozpkygspgaCHlW+u0QjsmHxXLChOAH2JaGwCu
yA9eEYGxtAZ9kw0SN0YKDmFZIVXeNrD6sSwauSHsorJnJP/dpHY8jIzq3GV+DvtqWSMzTZRPfT9A
e2vwYtjiV8cFwFhqgKgMXqZzIrCHSwN0DYKkWeDmjff+LZ3RtOld17C0Q5tKI+MBuE2/3r0GD6Xf
yQPM6XhNZTHC/0QC0GYwIxQJIYrYsCpojVFEGtG4+iFdKgG22+ublPQQMNhTV/h9eObQvElCj8/H
5wCC+F2cEAzTD8eoAhDMNkv6WHsysrP0Sc+olrei13NPvx2G0ZfkmaLEo1mRj4DQWUb83TIOLDBO
pknlX56CIXBBjjWAaR3FA+XfW+DzWM8ln36OHJBLVsS8VO+Lgy8NUOKRDgkz/S+GQNXhLLwbmwWg
qCa7wd5a/y/6YxbrWmhZVt5VSA3frRwCNeUJN+A2iYUEiH5BZFcoA48nk4Zqw/ZI6k4c/Vjpoqws
XzV2rWNBubf8zNR2vAAf7GIJv/xzM+GctgqVCV/0m45uEtxQmIcVz7LEf27Q032Zs5M/bBr5VnTI
qZqui7Yn/+iz7p85eT76X13d2NJxyskYdb0qj1Cgp1SuDk5+xBAgziZV9g2RsmRAvqGYGClaCywl
1yM3dxWVaPgaCidnlCeZ3GxuVFWZme4DAszKDAHXn7qYv+Vw7eKhycsrSegqca/KtJS5m1NsLO24
ywwGuW31zB5BoV9GaoVOOmwUedyFWRP4jn4t10oBvUGOVne5t9H1JxeGRftkVmtb9EH5oc/978Xr
9qfoqPdNgA3fEm8wRfRr5Blp8pB3ERNsqjcFPf5bszKqE1Ns64p6Di+U3NZwp6mADATpIjp0ID1T
S0wJ0YOw0Zso61VCeTS+C6qvyZssC127L9ZQ2bIc/nHjv3ITuoA6K3wOZKQncx2aeeE0Zw133haS
H73YhNGN0LfC93RBh+erIxGtnIuwiWIKOSj6BUEoyQKpGsVFKO8YBSaDFtPqcaRQqM1vt+EIW1/4
osVY/yKbwMkA06vqHM0inPK6gYTkh0A/axbWDT3/oIv0UezVY/BHLbtk9Eb3Vk3U3xjAVKNRFDmQ
ADlE3weV9vhAD14RwUwBSZp+niVnUhKlN7U9RSOEV8pdSd7zACaiIb0mYZEPjp3ZsvcyF5EZO8Bj
5INDZQO1J4AUL3RQoqjro0ckm3CH8bODnyd/1PdlBfY9LRA+5AglTAlucFjUS6p3Js0ytxzlEgEX
cSt24aKrv0TSGVLqqHzB3V356AKcpbZIsFrhUMIJOY/0bLFIXIf+801kkumQAZ7iQMCUc8z1huDO
rw17LigtQqajIYPEuQwujNUR3ce6P9qZdxXCgtWYkYHrJsIOf5JUi3Sc2KRKDvaO9HUZY4i+6SQa
4P36uZUBo0QEefIZjnEZNAcAFJkrUEQBX8K+LEPrXbm0krdBds0HwE3yahlfY2/LLCq24KTlhzBm
7/9vBOzf8tdMUhSiWwI8ggfDclesNuLYEBMQiIFmoTeBfgUVsGP3JumB9/0YBRXmfUuKX7OpKSmV
s267o/7WKC3QOnx00v5NTyasUH7kiQH5c/vi5HRHwN/mYm4rPoGOpcVPUiNZc0ZLLsSKhclcCIVM
NA/xgWJyqwt/bSR8HiG6o2wzotPaweAZ7oJAY06DblR6WheEzb3kfYPy9M7L6rMY33rjP2kPrnI/
lv8AvaVzszahoEmthKX1QUPqHmuGxTaLFi8sKZssi1tr7NuROWj0GKWb+HQyPAZW2U3bCTpWqgmV
xkekHsI9/w0DXpdHa2KCsxvhcbo/QpIBHZCTzrbQBmnH5jSpH7ySY34b8txwj7QfEu69x79aTZqS
If2V+47fx/3KCaU+PMvhIsMAnPXunxrgx6CSJ+Drva4Cucm5BFPTkgRctbNnAdtKADL8EmobTNnj
Hr0NPLY6B2iFW1xXgf5XEsZXe+OO3lCjF4TW30qju/1fcKeczl5GOT1PWmZqFsgguCWHCeKOKN0R
0XcSQuW/DcA7H1vAvG8Dl/tb48ALzrbNnNNwe0thPndvGPWkMBH2o+TcTl3hZoB4zeNBseX+qIXW
8/17c7H3NTVrfqwLypfpL59JyhJ7nZ/YWAZxTCj0tDoS5T923u8xZdqgJNEUQCGTFhxcjl5NiXj/
LMUJhnsbKO/eDQXMwNf3BDf8M719QoGNeTCZWLMH3WiD9yfsVbybg09iA399EnKVHaP6543nPVJ5
fvD0F79N02TPZ+1BRCJKRKvtw7BBtDcSZY3SCwYMOG3thHCTafoBJPPNWfHS/cRwF3ns8BpXhEmk
QLGogYgP5YVsDKayhQkAuhBokCiBxqta3DJTYbKamEoGdHJXjGLkUQM5EiHJXG7dcgESnklRaQKG
aX1SZXQIwmSRLMKHeAjSB4b5JlbqdWk+OgDx6MxOnx1uPE76Eo8LWAXOABjBHiIHi+9phtjwt+9k
DwvrZTDMMjFWH7YIIasjUsYej+t/WsD8LciTRhbal1DLS6zRsbdN77e2ap9U0Eku+MX6qlXd6lH9
sRJ9+iauHSmQyVjIYKHkLXpzpxVfu7lixaE6UpoeKtYO/7XAjmtlzh/3YRdUZn/VUr63y2iXR7m2
UmZrFr9XKhnH2uqgnEG+EaaeguFo1HPIDmgxbEI7z1by67as0tQLFCLwrnYnuxYgpsn+8KioQUc1
8BUKhHRR7Ta4XUv0Iv58lSvl+B8SJg3y0gDQcHEnZlOP6v/XQ7nUwyXhODJp7cc7lU3WUdSvy4+B
Ql6WlNrKAVv+12shTEWNnp2ZtqFQI4m8j/SjJSO6WSnFd8gDsplTMFtvFVaphYrJrTTcuqBJA9B+
2KL+6azmrmWxVkK3wnfMIq4LVIiFtab3MwZjXbWpGb/7gWEzjwuqnwpr6cufP6PLTAvj3looBfVB
0ui2rdkXhYVkYTWYWXx2pPvYNyRSDVs3hyk+uDMrjFRaXcl3XkjRCF19AbHvJLAgb1ov0H9qv95P
YD+Hy2kc09I/m/FMe9Uz4lJtsgr3ESXrLl0L1JjbQyyxhMKox3KMtzaPkRW9loolY/wBt13MG5pq
MQuU1IjqeqHB6jqLHiTen8CYxhdfW8tDYLRu2F6AQCDLAcrS+GVhrMAkWZ7I4UYq7NAdujdnPlV8
JFRHHO1nCfWQyJ/XvzpaeNsH8jS4YL4TyKD6jP8kGKY8ugt4BjMzweFBdxuwWw4q+pjak3GlF+cP
3w5qDWzxlPsLcyj+NPF9w8WnWupPKHyOUnEVE9PenRqMnYnB0BaPUHSUTH3rqjpVyCe0WshCqCY7
wR7vB4wsTtjywzEl9ZvttswEKpSyA+rvsbTFb2Wmc+bAfFaYJxw+QPxkD6vwhBFbWEsJ+v0cewRF
KqnWCHXQDSrOnEYEwcUPmG9UyvJDvGptJBYUHjY44WlSxYYasINcQv5GCbvacl2Ymm57whO5JhvW
nvk9pv/jAkpwq4Aaq1T9lmtEczPRy/RyScpqGiXk0yCSeTA4hmX2H8Oeo5mXK6yzKOQZBbEr3ixp
OHKWk1tNfd1Pp6OCXDinzd1OeO3m0Hv+1VmeujWjznOErIndyjnrcsK2GD4gumgGYrcHyF2iRB5/
aY9a+PppfjaxRoPF0iJl1QJI5jan2+yS43+UnMDDAaqGI9SRFgwqEwF9ZcapK19NfzDKqyynsr4K
v6BL72ISNa0iLkhdaH9gG/x32CHvyOe/XPj/apEhRqwaJJXK9cf3SXpCo3bgkkcNG63+yywMZjXU
6QzqwzPehktnRu1WU4iA4jTeCpqVWJr++aq20m+sDMLQjBcOF+NiCvjTqF74NjlU58RKzm2tcPG/
k+4x3R3EbtDUST2FiLcIH+eCMfg4NSWincdoN+WQfmSji7sSbwYCQBuVa8AvjpIPYBDSpxY8UM12
+ivLyl86U3l8aPLQcPzD+2IRt9d7LgIhg5BIOwx9/BlhJpSaiBK0btE7ILgqpaCJCFsV/i54SA0L
zo7PGyr0pFyBRv0VoyfxaLjEsHRhM7EcRq13Ac5JyPInfUGWgEvLQD57lu/UkEcc+wXDlUKsgomX
Zzfe9lHFzB+B+atsv1vPf+uIbksa1eWzepilO+a6xF2ZViIrf2AnEJwbCMGRBujnGalcy+HgP7SB
UIKUExZwE+1a/t5i5PkgB2CnFQhU83pYhewPN+89RRgc+ZorWcR2xSgvLI6FdWsUmXt3aPNnaly6
ZW//qsyKrNnKLV4uKRuV6248wCBYSNg00mKOBMYTpqHyJqHK89GA9FVRhyw9JZiAt6NjFCeTyEuS
o+MzmQWA7k5XYLB2w4bLC6PVfdNiCLLPO4nA7TApw3rX1IxzYWSo4/0X6NidJKFPkDuMVbNRJBdd
eFn8jzf3E8X7fO2ZOLN+NW+YQQrTEQwjM0Zs+N+UcSLDfuALO/SqJT+uq3TCmpU5XHniU2IRbQWA
dCFe21j4m/JA6PCjaQFt5Yy0Qcjjg95kzFYazf8GVuLeluLyOLhQa5o4HACFm/loSAsKM7AgZISU
qoZdGbn6Zb4VQ/HAliO9kbPMUvaVa09P+rKoqZ91hFjo6UnmxDqMODtoweD/5GEuHtbh5fFYz3YP
2qT93B03eFJhXUfJ748XxNFXfEknsfYg8FeGMYz9TrL/Utk5vGR+i+81+qWUIxiO4xL3SRcL6TPj
6kmzs9ynheVz98Bfg+hTbPj8QWRCdY5Ku1KXG7WUPXdWODtsLguT03wakGXh6HuuzgRCIfk6G/KZ
SK69t8JIvhPwVYLmLCgZkUSQ57bCEIFjGLly91yCYK1ndMebtjbZX2nhokDGukfpINIJpIR92O31
k6/m4hnrPOY0rEumtBwXYtO7jQCm9IBoPsozMy0UpVtOM86XMBfO+lTfkcQCPjtocGOYDQ2QSJfj
ea2GEsPMIAYp0BPTH1PMLaf2P2RtsMmyH6U5XZI1Lk5ZU49S8Ia76pRuHez7Ju85u1UUgJnvfahI
gkeCbdfOBkJxvjicdcRozjbiHxykFlU5lUw8uXhzff/gSoyPaTG26pitBx4d2Pb32mq94nHcLKw7
Ll5UWh9HNz46Ci1CMJpg+g/Nry2reZ1c0i22YFKKiCv00eoufIehXFt2gtf2VkUajVZkVlCVy/3a
7Zm9hVJ1ijzv2wfbON2hIg5oRCOwoG+ttzU6W1wB6lK464bs/jIZXwW2932UKPj8zUh6RbZ6J/d6
qkyoaFhUjD+CPZ7P1BrIdXR9do7hOsQyjM9AaOOU4E2+12G9SCu3yUftpJYrwjfQ+POffk+Bidjc
0XY/75WgwSndlmlPP4T+5/epvkDuHQKvPBrmDOGTcapHS03gQdL8x9FGSHXqvkSib7HAcsnSe2y3
pQMtdI01Yo6fYRk+OKmN+LuD4lFfHfbCKMkSZpxG1yI4hyy6UqTT/juvqX9W7KrvYIVUxblb5BmJ
tCmsSG5P6lNXFUwUZeTQgfylZMUExnQczupbvSIRxzNjA/cVxSB1SGhXPJycKRwr5IH/aihK5Wqo
Om/PeIq2BdxavuFAZQ5vNg/i4vkZv7r4bkA0vMWsdqx6OZMLzELbR78X6GDgbuYlItnq3tCLz4vY
Dvp44fSgOKuDAu6yhBKimi1iown1rCzyD8OWjrYaaJ7vEl7WCIkqAg91THSgcVEGhBQhHJn7sbKO
eayw41KI7/7cKab+GcMBKZqoDTXEMoRpMQQobmG8Zgeefi3G9Z5L40u6ZXO411+KXB+4j5uqHbJZ
67sz2kSbx6i6932J9gJpvtSwFfw3kNbUdnpM+Br+BQitquaI4Py1QS1znYnHDeMOw62teNlFeH1Z
xLzC9xeoz4Gi3x09h9HEQHWLKUkQYgU/i/BOG7ihIr0/t/0SJJj7FijZ/nSXW0fJkAjoY0G/ohYE
keqj5uOiIgCd3a4UzyeUgynRJiRitsz+CVrN+oyid2AFcBtyB7qBlfzr18OtfnmviImG64rLWroh
Fvfrx8MWZK9ovNUobi5ymTr4P9ZPcA5tpaYzwAQMbKoO7J/p3aARysu37/BhJIukhPPra520jk4S
+597AhDY3PMUAcFUe5aVNa19VFctBsiNGk6ugrTkKSkRYiy8T7ZhAf6FxAjb+/+WlJiGZHTu1IlW
yRzaYCPKENBYJrOdC/pqdQDTL037rpxW7kIKFfWHp2bceF+9+hUp5a8tDqGV7MT2VyM3OYzQgySf
kTmo7a+2tBKBOmtuWsGVqjZW2VpccbpJW2fg/tfFs6OHylxSGRA/Loxw2pAV+CQA2mwwcNNwXBSb
0yVH/Lus+Q0KRbGW2niXb1DRfhvp8V4U6tq33BgcGZQsZCVGJ/PCXUukYIihe1JcrTB2TyHi8MaL
e7JBwD11p2VXGHS8C6KGqrjddjhRSmT4fksyIVWOlVHPVH9kgXpx4SuI8AYXIHL3T05STnxn47Pw
BD+am06v990qDOfZnDzKnx8StPnFo0ihpjWcWr+rfPXTZp0Qb5eiZY9qOzO3ckKimAGZuisdA32G
qJKGclgN5rtPUnNUo7g5bqib6J0hDke77YtG8aJ3/NdqUNBFt72NVNzflpiSAxM0B4y8Stye0AEM
Sxqso9ni9whq/p/NhtuSUR6sABno8jSBZ3VsNU9dPJdiLe3M5nyH2lxH7Xv49HTbCLOl3h5i7PvC
TSiuOX+HQPUBRBDmbzGTrfFfpE9YeC51W5ORCFkowWm6D9Bo2pU174nSvDJJiNSvpxr2AVXEWJM6
pUGPqnLvUipJankg/c6iXr96gFKh5EF2CpZ7gq+22bO05/A7QhCu2QgjU03VS2mDm1y8s7sbZQ48
SkdDGF6iBJBjAQOR3K7wMzhWcZxex0JemxIQNp7RFtHVSL6flXLz5Vh/aT7q0jt2BmEpHnnzGcyF
jy+GYJgs+wZKXiwj9yejDayFW8yrzuNDYY76SG5A9bRsSHIv/09tjkeo/ez3eHQxNUk7WmWs9xXk
VKLXgx/998I3KbSKUWrQP/+Gj467eGl3vJAzUjPM5gE3QPrc5VtMVnQNnkRQqWBt69nOxv8oQzyJ
Ve8YvLU1RI3S/AuxQppGFitLmYi2dU3nl7VYn6cnr8nuw1He2rZ8Kp6LoJdWyN/Jf22eUdkrxMn8
NfurZ95jb1C+6DNJIdnXQQD8LNZTHzEywPSi73YHe+wy5ujPA4y7ER6Akw6VMQ4nM2xqhXGxA8MN
xLam92ahxERd/PCHQ0DpVAOYwraxpLxaCXzPcRLv2EFUzZ5KaOowI/amK2h/m6G1pSUfMAk0r19m
2xJL2/Vo6GdCkjvVqOnbUhfvKUqa87yn9CT+KKzGODOR5qeQsxC/upfn7ccHIpoezlrOby18zzWO
ouotMquUo9l06VY6gTFoq5hova80SU8ft9XikgqXwQ8lJrTkhP97kJK91dpFkVsWnHSOLQBTqyTl
SZhze+crk0IpFRJdUZGNrBu6Ms1Ru7MCSFRvENuDLn0nEE7d857DLqaBAqXlVocZobzeTMj+RV0l
BGIkuE6LOLdYb5KmmJsF3/apcuxmcUxyByzODkLEBWabV0iG+gMRM3kahTUC+7Sbcj1G6baGmDlz
H7LSrR4W6WZWB+C/4r71CNRn74UpF1Lb5jw37tEWhxT50ciiVhN/7M4hNmp0duwhvPzH3YsygBJC
bKlwu1KhMQqSD/m97MDyvoMh7qjlLv7cOxbwDgMTml/u/qtjcfFtyuUrSrWtHBllZdTrKTjI9gYj
j3W03ODCGP64vEoE+Q764ujl7JMp6cXq0Aue5i1TngTbGTIXnyOiID7w6QLJM5Irw0PObpoePcJV
LqJ7pfrpIuTzxyiihSc3XXzRfGFvoonaXHn0vZBrfWjI/dNZ5q1/9ZKCE0/lptExjJTyYhUGVPgE
6giLwpCqccYNhHVp+3k9+hTgkpkfcVtvl5FYt9fMgX8GLAfmLJhJEaxWbEv2SsLPjThZd0FxlVqo
bIVvGjhswmsbPbEqNlRRLQsXc5aHZfmfjYLFWGaWLEqWjbay94c4mtEg0FlL3KnQiJtVE7esmlEP
OtLWHL7Y3Yrl/rKo7c1V7lTWk/wGhMtXjihJ4y7IyYKosri1JWopA/xG7eNjJGPeK3oaN2dHjAie
vw9DW83D3eJCOyn5Yq0A7ZD5jNXPsA3eltG7mEPKWRI64S20DgWgZ7ZcFm+F7uw8JA+yu5b+WGcC
ERq81U1S9tPmqlgA64YI3BhLqwGviL8f0QxLIGvHWWCIJkNWjDeyGOyo8dQFBbVy1YeBoFOm1BYR
tU6RoldmDF312NqrVHPuP9amHra6GZeK4XUGyNHU3Daqus3KvCEPB0LPNF/NBr7ZdZ+JoDpSSdA/
p2AW+H2Yeypzuch6GQsTS7UJBaNjtntSbWdIMtN1eBUT67CRtJO3bkjwgMOFynyNBsdO6AjnEMro
UcgAqrqDV0EvyeDheSf/x6o6/m76rYbe+YMNBG4rG2Y8x/Vhd/BQ/W2VJiPAd336/IXKVpHkaOtk
lV6xdEfnDJPimFGorDsLQpLQ5wFQWEDAAPSQHwmzCthffyqFayDs10DZXhY8yltGIb5hoHDcRNOj
g3ZlBYs3UsX8fkBHbemgBle7w2MDpSMmCoEXkgHJIGsEv4la4ZzA/O5AULKBwxe2kKH8qwUqKuc5
8D+zlLfMGcHYOs8pFQsKWZ0YDpez/f8XfZXeURdihNLPwE5HiILBFE5J8YVJrFU67wqQ120PjP5u
A1UvHjpZTP6FZpZzFvTt2SgRCgFYTUI2jJq66SGw76V1VSK2VavcBc7e9nyLDZfOf5d3gGPHy/wA
dPwkU2PAN2q2OGLMarXc2dJA+oHl0rFp4N3XlJ5510IqPupQjMkACC9oLLx3ozNsqArNF3qC+3yE
jo99Y3S3gpexbpUk652Mg8nLdYNP1cA7k4nRcQqNOhwfPde+ed+pA+ArGX01kUFyi/RSCCskv93t
1mHqMwvtUwbxkGXcSG1FO1AYZRjWXRUT52GPKPF9DeVugbEcF0EmeZIhQdFmQ75CSrHJ/5o5U29M
E/Dr1Y6JQgKk3b6Sn1djzoAossUgomjVw5U7qcjSJrHGtoGaNoCAOj0Nhg8hh+juQ78hQq3god1v
GEDW79XUooA+vBfQgvqHsHkC8GoD99AtN+mQhQb4Qghbg7ZUFEUw8G1NrxF+W97gLb2AMZHVz/lN
A6ULiDSvpT+TVqUmZAyO4k6KEdhgw2p3GTcmdDFM1Zs3LBGGrjuBF+3GwDhbEUPP5skt4LsrE9Ra
cwgk840H4f6gOo8WiX8LT6HoeEGLEDIap5vv7Q+/yFidSNltiPgaUZE7N/46FukFRlKQjEQoaF30
JS5orLbvy2+l3xPKMp+kQrLRZGvG/91eqcl/QkyAYTuc2nmwMoDNFwf+WuiX5JSFyiMcyagAlGZc
0QKTmrM7vR7wxsNeQahFi/7CFX+Iq/RNoL2ErGgmWFJB0Fc0KPh8sylH4KYRrb4slu6o6ZtvDbX1
j/PQvFlQnxS1BPF9tX7UpZVeClBwEvZCxfG8jBgNSgelKoZvP0EeRmhYLvU/UKTdHYjL2mwUgZM4
pNuOp/YzlL0XV/g//JfqZevA80Xsuy6AqFsaJ+Xez5KvSHoKlV7YQml6NrXw1ps4+IXMLALLkrMe
MZYObOEIJ91LQ9h3N0EqRslou6rTY7CQekG8fZRvo+vwUd8b4l2gdb4APPgag8tCF+wikeuSzJ6N
7dY7sYhzdkmVgO1k01LuEGwpREGR/gs46yKGNTfxVQ84xVb8CJhhQFT8vEbwnUU2gX1G7tPDXCRp
iNHB+HCu/8vRJrsb1G0a8ODlMfxdSQoPi6xEqSIhRjcNHBueCDA6+81PadNK/BEwSTHNGKkT1Dw3
UrOrzM8hj8p79Fa3ODcVlue8Y9hiWlgmHS0hP7+Oh22KNVYl+ecVmqjIrn7LgVy+g90ab7aWVcEb
jsqGj5mVNaJljmLDKNOtVL7A4eEQsAMBilrEguagJa1XwEEIv1vII7PoXb6DSdVTXPhPf22oh2Uf
tRdxdBd+EVgHVmwbrjGG1UrLeJ49XnvfEmsGs7H8hMy0slGXgUSVZ9NCX2P03hEVqwSZF13tfFTD
+HYPu/+jIhCCzhaYQCnieV666ZC6dFmO5mIrtLufNVIFL8q3V6qWubVojuSiKyrc86PeXTpR85Mo
g1XQkrUAHrtqUEYrVXHtG8INbjFNloSpDN0XK3+v42kGD1tEWITeEgBDU4OSXbZnaUkWsUSPCJ6K
Tq8Y4BIx0DzUleH4I3e5g9DFIt7QVPA7h/oT1Z4SZK2i9Sf31F3oZgOktnHRTKkbnb70otQTZjrQ
oAIdpYW2nTL0wujACXv4La7TgNkBOlIY0+GqW/yn1gtuOczQIDn3zmNGo2kPJ7V7Xnfp2bPTHfrP
fbuP+AK2A+8X6TA/vMrpw0A70wUUq/x0eXbwRGUeEi4f7gq7Xm7NWwKKT8Wl/i6g1CoNieFNns1O
ppFqucnU0D1EhbyGh4brVgfBUUf4AURRwtB5SGsFfa5WqjbR9QSBpnF0M+NkUuYs7y+wga1iKQN7
puJ2lQJFmPUGGrlSFYyWBLCiJy/bO172Fasfa0rxnO4IwHkshrzA6g/qO6qaZNgGdfuqC2WVCva8
T4ybJ2IBjJXuXu2jGmsojqjxi3/35Vsa9V+YB0dpEP6g/BpnlXCDP5gQ2YQx3N0q+mJW3ZGa08IK
G/Wtz7HfXfZxog7zjGlwX4A29rGCzkbVv/Asxr+jQ0VZ6PNbpxVeA0BQbpHzxJyHOd0Nu22VL3d8
oMrqGPHuVmS+zaz0pxnnkWQYtUAhDu1S1XnFkl9HaB7fKd7LRPjwuBlK5RY/qtpqeFpox549hX1I
D2v6KDAj5Qpy+FiHmtC2/plPcvodNsDN9p/RPwynsrz1jUbDD6kNp5xDvKbbPJDOodnZ8rVn4wBc
/r7WjW8zO1EnaQvS+29Oz5Uz9w1gLtba0ai0ghMnwli+uoPBGwYhUzDReee00k5GkwkBVm84+l5X
YMZemEa/srYryzcA2R4rcQt2rquJ+IF7wvpnOQnXNGU2eGm6S97PgPYxLtEe+q1QKih4bNyXf32G
H2NxRC5gxafSOu5bV/P1KdYELCYSHiBRwZ5fkNX9n6G4oZIZpv27qeSlZ0tgFeqQlRwVhniKVEwU
DwWdP4J83/DETh6ZFr9Z/bTjNzs7YLpLPZkMmyaFYA/7LL+c5OyAky1G+8iKCrw5OhbjEA25j1Fm
JFqR7PcP7+lqAAyR90TltNZF7LFqZUEwPfDTZMbXi40+XvU9YgPbZcJytpPkTdE98UKgeEwI9Wrj
NkcbwGlmSNLj4zT9MCl6H+peTqSi+8ohs9K8N1AJVmWTK82em0+J0HrU1A0MgbM8GsQRXgcIvRM1
xkWfClWkazQoxzzfnSQKjKGdpADqIXbkmkuxWLGTrqZZDVHbKhXnkwOHOk1lMaqkKJVmChCv7kVA
gKwhG1N8SQtotLOBmWqIzfu8OwDpx0Sda2LwpFnjuHM+KokwLVqj47EkUDJjM9ecZ00BZ2AvrjHb
lhG8I+vN/63Zt8dNGgeO/MmZv2tLZ/Q9aL9KvqeX3YH+OTtV7Jj06DjcEE8djtVVnOChUJECV+FN
aIprsHTdQROqsu6dbzg9G94HCX7EdZBXqd9PT6C8DDkjwagWJavSP/qDOueZnrzoEiQpZSVtCB7S
uWsiFXFtlyUUCaz1q2V3WfbsrJKwOXg6k2BVC3S/ZRJ7jTCnMzGFDN7f1VSO66b12i3p+JS9bABJ
IPT+Wsvid5Gusp8rb4N/IO9ZF2Nf0aRY247/gNq/WRZeDRzQo1lJfg0GQc7XEE+ty2a8BAykknXf
3DylQn7EpH3uiFQ27WOYz+JqD0cvtQb3CyLOARrykTmjap2+IV8zJ+kWblQ5Tn2rXXD1g8/OLLhN
0elUZl0+tXjKLm4Sw3Qhg5sNlxm8urHSdv385iuNrBKX9EDdLNoiA0fklpgqtPf2FzqRJX9AjNjZ
sF4VkoNIFDQbDkv2EJG0pLivYdE394+8nBiwY6z86W8NkaMIr4EOz7n7KZR7/df1BuqbhXonkQro
1/eqsgtsK3BTG8DhWZ0z8c8H0G4fqDE2SlwNMAzPDFeE5KYbhYh4e2uRAhVq0kmayoi4VuhFdD8p
91rs+UUhZj4srFJU3CzpchEGkA4D3YVW3VVgGpujaM3LqreZWgl4atHlOeOAxYhyCTSaJhXJLM/t
mLyDQ4OkJ+DVqUtkzqM0i3WSy2L/I2MRd1FlAe4LVEkzGuWKFyO1nNYyb77CjkKo5Wwh3fQIck98
39QxQYJjPxE+Y+YJab/+3RG0oQiHp4eiSkOlR3fbgp+c3wp37iohghEsgHzQO9bWx+XaMNVSHtJ4
rGXI06VnoKEGBZgRd6csdxIOmOwNt/exLtk3fDQ3QZzDviNX33vj1r6uUm6HbQPUs202AfSaHvvp
4qrJuEUoEzzHYXoZ3/yThnJkUslW4To8Yp7Gm+udCKt17UMDqv41j6u4gqf6e+0ICSgc8LJjwV5z
oyUGPJfwPKmzVqZ7Lhr1PHKEEnsQyR/miU3VvdgEc29H0v+s8cJpLWDqpvpJOFheK5SsGGy6pC6+
x+fM2n2TpiOAx//3yvJ5Jw84+FGWQS/SoMm2X0DftfdLP5HeQFaoFS+lfY3rXUKOahcER2rzPkBU
19hAWIub/AmKho32/z4xuWh6/9DTTThnSx9Ph+RA6tU7a73s0ALaHNsZIKdPIodKrEloQk7ZRR5K
sk/ocsV1WYOrmbH/wb1sEvxqV6ZdbQjsUJxZtXzli7JR6wP+ywvERtSJHgpz7b4/YtiPdbt8zn6j
+p/5ieBC7SFZnLi7ukq8i1q3c3stWr7zRwG/8T5CE3KwFHRxAyWyGbFpqbiOWqD0y4WNT1CLEn9v
eO1emZYa43dllgiSnMUKJ2QWwYkO+OOpZmJNd6e7m2OOnndhNA+xWIrNY9lqibU0a3+suywO/feg
/Oj3tXnrkqBnytdq/Jwe8+bLE2tD/CExUUaTPIHdEB23ZAhjU95qtZouh5QUeww1GOiMQujA3S+u
nVPavQyzcU/pc5/YLa9KC3yqU0TL04wazDF1MojiO0+ROJwCo3iv8/uwL9Smcloe0MPfMHj1QdIn
kMf3yykTRfqHVY7WF/BpM/Ny2pxRCM7ayXnh11qkr8jLhDyBKMCyMudjGwVqwOLZf5brg9c4zQVJ
zag4fL5XzYbf+eVbMoGYDEzy1/g1zBNHPiuoI1SCqZf5lfCBnJwD3qQ5OyfBerurM9sLuKZ+7LS8
aOWwHtDppaNn5gNTelkjW11IrgFyG0QUTMPTMuRT5UAfqqv2NTLsbHhc9HYwzIZATuLsTNWmbt3I
7Qsw6fUu4ikt0jBGqKhVGVth1ZBNanwA0cYmNXII/eXlMpQdD/SIZyy4dXUT0H9B/XHHMgQdeor9
AfaLsGFCJjc7i1QjHR1I3kCdfQPrurWGeBPwligZ0oCA10zxk+FL7AOITozVQVkuT8/YmJPM/WCZ
Y56jfXWJ5lYGNXb0tdc9AnSn5MBdi4rx3ycljhR8kJAjYBzigPkOHgzfSjuf2qDATsxJsG3wMZnw
noKUQa+qid3++H/8KIkyjiMNwquRYX0sVA4JTShGJ71+BKoKk5Hup8XKi1k4fHhpCXf+wIthdbhu
S+dgTb74qQ5YP2P3ETvYwl+vnl3pbmnpnkwq9u1GQ+GwcKqX8eDMDq90XzrrkzQ1YFbOU0vccHMj
+Fpu6nZvYXngRFok0f3JmSuz/qdSDYBkkBrwo7xcbAI4sehoXfbBOk4k7jeDmJZM4+It+Ff7r93t
sOT/Ezlo7uccSRB916W+JjzMMyJ6D1Dq/YFiwOi0RfC3AVZEMSQycOXmzduqUUtQATf0FTvc8L0S
93tt+18vL+6zPZmo8obXi+pwd78FRxRSbN95s2WlQU7z+ykQxpHlXMkUmEBj5PeI+1/lFywjaTFi
kdNfIM7FnvmSPgisDKy1TCHsPdR73wTzEZKLcoMvfjGDlgjvcSBF2ybvTOf3EWcKOw9DaDrCHpGi
4thBFXGYsuVe8EznMKmJjtiAfMkiUhksgjvobSQ5V+d6xk1O4BmGKuszlDGpaQ15JQ8G1vACYTjn
i7TVqyTDvTe0uMf/X3qlq7fpOM2Put9w99grcjrI4xrqgMSl72Fay3XWBukqE/XjL4MbhLeSMeSO
UMsw0omwei5skKQwQi0r/Ay1wecKK70v4oG438vqBB4VArEls3uwbVTScGK5a3B1j2kqQ6IaTl7o
hBlGp/1AfDi6AgYwhO2sRyeF28Hc4XA00bRUSUlqrOZQfW7qaSQCb/IrtiQzRMmcEchAEuANRxUh
uRgn2+mMhKl+P272lq6AgwMEWt4obNtHxpw4cBMhGIECUTIxcWXodpKxoTVPZkHP93u0u9xOjHWG
4Gqrudjz4j9oZfhZYc5jwN76oesg8b2i0WehQHnLi9yj2WXc2Oce1fx3cF93bW48MLG0U6Mqcmwb
1VwplzEPW11k2/FOgsnHl7N6wqInJnuyyNPc8YuzfxS6pZ8SSjpmNB67ngNNbjhjE9cucGu59nGb
+YvFE3oa6xo0OqTdDR2x77eeMbqnwSNmtJ54yUTXhBnvsKQkD2icunmwZBXl0g7Bj3AtmQRfGMeE
VG2MICBSP3hsrjxHkTUOugvf1DM0TNs39vBXDF2RoT7myqFxb2I2LAaWF9tihN1BZfIJDFn2ql2h
qRFRp48CiwDuJY/VHk2LiE+9B1WA4ozRw+8O+enq6fN+pBeIsF2UfXCSAPXDqv9pX0f3MXeXIj0U
EuRBAfug06h2QdPoOc8AnKOLsKx9iLt4OciBT6rwEhNbTMQViG9DR0AGXwj1CuqMpcyaM3wcm3vW
SYBYxPDcVJ4y5OAbdv03kCjlH9kzh67cIKt76wyIhoAvrPwZBkWxy+5zXBWp4uhbOyRmUJfUASmA
AQ+sg5tNCvVzVxCBr+8X4wxRr8YmauMlraK6wrwF8xLg+SVm+7k3s8rWLCCBW5yP+NsKukUhKbuB
3q6qd7CzyTRmz5XjzYPG6XcA9436wDl6kvnEyGaNBzx3B5nxwHKnV/MhKBIsFdypLNIITcgri6Eb
ov5xFRpCiWGbExVJDDSZZXI0xFAf7eg0mjl6i4wi66Gse3I3dvgvShEy3WdesPifIqicT9MnZmW6
Ba8liAYAwx41/LPJYyClZRXGn8vvV1AwjgsmYprhkgwYe9SwWKjhm7SmbQsD/7/ZFkWLz8+v4Mm6
OWzz5ftrmbM8HOjDuaPoj6qBBqrqxv8Xj7F5WUmE2WOfupc3SuBSCeMFPwjTc2fMULJ9ax3Alvdy
BtoJpoP9bkhry12JJwSDsukCkw4yJxdObTcyV1ZBhLfKURq7ZVgS+uQsdM++h/W9jq0g8KmgU6ur
t/xJ36d7li2lD128Yq76Uvb5yQMzP1TQ5qyVDg6qk6dNXPDKKSwLTEA+HnRRNp6j4icj6LpqqCT5
L7Iretzxm/bVuSMTavyCe3wqYUTWmQkuGPXIo+J9xvN4kUAm80fOqO2Pw1olmEbflzdxLyL/GiIk
XIJolsYu+tSDNPZXE++VDdFFEvSicDzVPOmIrq0RETub1IDoleFF1NvoqFZLGc5vjsMZVlsD3XoA
jwi1V30h137/6g14PERvJ+waK0tTqzhmClaPZXfKntyoXmV3pIi3I5SCPrvIwOLjkUfXvuGkAFL9
P9v/K9Q+nbH2CB4BMhTqVKwgnR06QLeNN6MY4+qkoQHqJoIpYyEwKitrvWvqzeJvEO/lZYpFJoc2
9cYziIYOwlO9NSy8Hnsmz3F4ssi+I0+J4daGHADlZ2HB1wPs5xC722ZMKV0TAIRfqz3TQpsIwnyi
rDG5N8Aira+U2qm3noj6NhvBUhEpwV3d9vEZM4RJqkSp1633syEf74bi4C5AWPKEAwmlH21iP2TZ
cWzFF08SAh2d+WkD7ozwadLSsddpoPfl485jicntCELmwwr+Y7Tc+ErcscYZiMe1yb6rv1yw9uPG
W8sjLTDm8Pe4aLLnh/2MJnHpCXe4ycqOKDVcLcmKKAq/AmLntbdCsaRjOGRYmRb7GBWl0LTPbSfs
HwTCjU2mGXqZ/9QFcznni2qWpEA4G/0TV05E8wAZLz/KVPGf8UTT2ZXxx3WFBTzuRB6S8ZYgnv+f
237TRC/e4742Aq/m14yviDoXICMoj2IvJ9peu+R26lF2mNOgIN8Rsp5AX/Sh+/O4bsF9tMKE2cAS
MaOWAhExeJsx/oFciBbRykkqRDupoeAaa3ZigVu1XWWs2R2KWIOcn5dx0f2ukxsQsrZQO9/gqZ+X
Y9bVUOZCoevN/FATuZjnzN6fRrWAERHvHfEo+zSE9RvVTYbjN6IKAmALt6+sTSYla2PNGr8uVhZ3
LQOUCyibSuH2IfDaCcBMamuQxo3ogTYl9O5CM+i3JDz11Z1vRtZcOU3JyHcZ8bTHY7J9h5WhtiPh
1LBojExM9tP8REq7hHFMlSixNq9hScnzAnfRPiUmLBaaUDp+FgMHKl7uaTW48lMdDsS8tRqXCITh
mcAnUAoR9lVyOROtb7tQ7Bm+TsSjWfN/sU/9sYDe2IyzK9NrYUoETxBL41LNMYha4ZdWRRI04fJK
OwzohVPt/x2d9Co5zd9mhdUe7SMVn84eTfrqLsSgytvkYZd/8Pjxd31cbIzgVaO2rULioYFgBnRH
INhEej1bKovc2Bwt58hSQL+6SnQlou5kWKiME49Y9RLce/coP5iftlt0Vdt/224ZEh7xBVVcMaVQ
4pfSW/4t+50q1IB6gNW7EbaJR/8sdRtLrcbcU1NGEEwqB2hRLFtjLPzZurcLRWVEW3rZkzbogYHn
5eAfv7k970yP4uexIFcalwyH72w98EIgv04g9O6u7LVDVwAPb9m5Xdu4Ft8BKqDb7C2xGONwY0UQ
i0ifV5GpTCBrZf4r72VotzdjW56eyUbXtk6mAr8nMTBV9stcpIkc9jfV6G41FGluEAOBN7/DGFt/
s0HNySVAG/AZg058LSjO1WydCA8LRk5JO9LiUXbd+QcTEKdziso/ikZaHXnbXqFVWaUDJJPfnLhf
pYjyW8AhCI7o5sbvN7OmRRE4nF21oPF/WeUjy/ECdqqTJm2mUZajedm7IpId+zyhaMXnMmem11hY
JRWPxcIKe0OIy6SXq8l95cnDC1QdIc0mD7x+e0dXSDk7ZoUmydo6+Ppfp6+6ka5ALLV9+ZeT/Q9/
iNI/KTyCoo4cxrWa4EoK4/1MydKm2tqrkEP2/FzYCfMcdI/ih+T4z5T2gd3xRThb9EG8XIn+CpBF
fA2us27y9RGvSld1GJ+k5q3o0uUTBhtsgbBQesiXq3HvotUWLUGzdMi7pXkdhDblqqwjpv1rGrlE
qMPlgVxP9UoqsWaC6Rv1TzCPRIq97GQvsogWVXw12/IYFZfOUFSenMtEwhMnFU4dHS3Ylhw/vpUL
D28Cmz2DzzFKGYFaqWM6scDm8xf6Ku0gz5LZfdXQ2DGmbWglToidWoVWHXk+swOxcJsozhvRIhpW
A/OKEEtCsbQ48Tp86zzwFoefiXL4bcIubhu4DFRvYL1ty6Tu41MZi0F5edMdtU0DVMZvuf9UsHz5
dp0xU5njSSfgGAgWF4GMfQJ1MqPL1zuZYVY0blbQNg1DF8kxHxL2vYvhHjEvZJqk3x3mMbnQnKGy
coRefiJKoofBh60CHpT+fPk7vRJF8PcojksZUKCqiIevzwXMi0YimOZf+vbOZ/7nzE1I22UeAjcX
EICTsKtJf4GHz/OUW+NzpTSNQYSOPuWcmNEacSGPesUmMGPY/wL19kx9gNEbVYaVEYBWtiVycBqG
vtfK2fNv/5Bdn5HNOMyHfV4j99WNOtdjepZKVTB+k669nkRuZStu1ynGrR7sGQFaO/noiZiH4WN8
9A+mjEq2NMElHLVKygzr4Shz8lXT8KMmMWGaiRW6hcAcrcJpVhnVQ4pb2rxGvjjMt1uPsXkGUa/O
lESTp25ZiRwuNewsGLnQpaxEi1OAZfpA4SjdGvqX+Nvfmi6CsvUKbcpHOxE7NM3AXBsyrYal2/TE
GULeqCS9HM5NTLsv5ozgPfnGo6T+X1QDFwHtmsOunf5kgZk9RcB2F8DJi/Owzx5lRjq2q7gfBj13
UJ17D5tiP7/I6AkQYgCc9c6NIjp1mYzssiEiE9ITorFSyq9IiP+00loTJvAejNzpgYTa1DUgLYHW
8R5OkKY0gtMM/WnziCrpcHSYcqgu9vnLkGNqwMKOUZHO6IwdIu7PtgmN4Ghxhx39fQNRAIG/8cpr
fKJMHwHBTLlkLbc6244xbFn6OxxOlQ6Ge++X1WOPzhj683DsJaXH0KqQ7t1C42MAIpK8INU0lsZo
nwtAoQWzaEexS/eN2KMkB2O0gc6U0Tf6vJLH+ax7XcLLqNdVd13HC4eC+35hEqcAwYFcdOCT6M2z
3q3sbCXZz8GZ3rbAXMaiKovT6eBXUbvkFwkVTcS4+1TnmKQyigbcUNOHz2NZcGWC3nSL0PD06of7
bEqB08uZwT+/b7mYRVhlJjRVFatSMcEbjPy04w0gXyMI0KZQONaM8bmHfY4x3qV4rO9f+E5JSsPK
j693mhPzEQnCGyArBWUejSM2i8mtaTA2NOf027Osu/jZ2VTnfbXvTYmScg0IBqKFVXGX1rjlyAo8
qKgnlon+Qqmeo1RCL+n3orJ6BRN1nryLrSD4SHD8/H+ihfRl1u4TfM30XoJlZC6mo3l8VwOmTeU/
mSkRf2dofHPYWmHIZms+XRuVurmYkF06qV5TiFlTJvtPnPkrm5pqS9njA4+1iNK+1AQByyfLg/ss
PGkbe1j0Q9mmg/eYbIX5mySUdhO7g3PuRBFXvacW7uN1+pSbpnyJ1ovkECvkNJy4pvMEciv6fkH7
RQfmd3wyiaYijkK38WlW5DvY33wWvexa0c0AbqXTPm5L7eXZFrjTWJyc7aclil6y78e+gUKYFWyE
Ug9peMxO8SEB+2JArk3MQqGuHhujDS3U0IZQ+6Rz34yeMou1XNWJEefJBlX1Zaa0dDHLfg/0RjWO
deJBig1m2iPgagNhbZ9/5C2558AXNnX08LQ0OD3EKbhx3mhbAd060nbq+YJS84z5jrm6KyDw3dEy
HmeOdxoGMThx0Z4C30nCkddfoZQEdl3uu/jsOy9PKAXzYzVmcIwpuONomFcERPGyNoJ/9SPi1GSp
ZZcYWAHejD8+Ye7TcDz6sGJuvo0AkX+GnUdqHoTwLVFX1LVC5GceK6P0GNxWMp1KmiB7UCpSOMVR
LYTXH9ApZgMzQrIE7pkM1FaicAJHss13op/iL7+lmEUSQZ0cJrb6gNJG0jV/yRcGASfEZ9Nn0CO8
rUr2ASYDp59mX0vOCorWfut9T8Qi5hgnihdaA2CzYBtAYVUFZmKAs4jGn2ywQANb4GAW3Y4FG9ab
Ft3czf9TUypHTAGE0htQyM1swKREzHqBz6l7O9M+3p/kC+pbylkJ7Vvs8ND5Za9HqRbss7kqw/Kz
+0DarB18ItqTjZphkX4hzj4DG5Sd4h22DGtXFlNZIBpSdiCbugUU2UFSb2cWHZMV5WBcC4yVPHSS
MBTpYupN4ljKzyvc4Bxvr2SlIeq8MbZ4hTumou9EZhOHqyiqSBFEt8Fu+V4XsXlnxhdSFYQOi/Mz
tSePynRNFC+CITjZAD4V8ftv91h3bGruDhnXlJnbFJCnSIR/giThVKMRgTngwwakNml4pjTx59m4
HspOxj7jkXrjmagTPE/Fy9rm0YyF7C6v0K5JXvQQdwJ7kzLG3DXzpP+fhrJaTkKJoGeoa0atJhKy
Af6oKx91CYV/akJ2CDEiheJd76Y7KtALJxwLZHnjgRCOc1Acb+aYrbNzmFH2GRR4w7z57/WlVC+o
W1vapuwHARqTAX6QuZ8LdVAzwYu3gjc4/3HuTm6oaY7axZF2MSot+bWWElOH8frAvB5r/JYQmnHs
qWs0Z+x8TOKACh/xDCEIaS71IaxzzeHyidgY/jIwsQZIoukX6tyA1zkEMknehnUcR+32h+JG61pH
e9JGieuJBZrS2lcqk4q+yoP3l2yxbMIsw1tbOYpdMRqj4l/+Rr1xgHTiYycUshvB9CdrxqBiKJW9
25BO4oJ0kjWKVHndoyDNT9SqbcPFdX2SM74iquFdjN99/ykKZOGaim+53wiY4clSj7NxI0VtLkPg
PntT/c2K8sJePfHsK2muYKpAxZ1tZ6FDaCT0rWQ5TySHJZzbM2ottyAZJXSmX94rKy0TcGb7fv+m
7rNScwzam4ByZ9Zgro890LXx7UZCNQ0932qoWAfEkA5xEKmHv2SlHXIVwY/BC3GH/typpS7FfAFL
C0a1xvkQ3s03FggTOpWc66cdJczjapnc+9kN/xaxuoR3Loqj8HXJ5Kns5A8jLEtZVbfJKcpqV62O
WKf4FTCVdDxaJ4uI4BxXwkzXfZJbfoNVNlnHbZRkusmuH5gyHuBDx7+ELCyDyIcNQuAFAF+WEo8R
6RQtv25vULLZU82gcHx3Uz0BoVNM3TNyZNTf2DQRsiGSfe1h5hwrU72It3ueQikt7fBvHvwX0D99
YUQQFwHmhwKK3/uYVqY42y3yfiQgqL7JFT+kJZCuHLv8py+cZoJH7YeQ470WnSQ8MszfKHFPuhFO
bZIZEm2i9fUgJawSabIwK+63M3dPH5xUqH1MjjFQI0sWAEo6L9KpauVWWqsZr6bIQ2t/zrr4gxGH
LpRpNRsYAjh02/qMM0ImMZJHGijAI9lp3/syHokdJMd13E7XWvUCkHrRaLBHaLjDxKufD5uoWK4C
NFlps4XicNMrakAgC7caLDyonRoPBEmvUolr27IxXIbzRvun4+WC2l7JDD/8PNqnDrOCZtFPIoYo
F2z+qkVpSGM4VKf14eH8gkq5grJJrFC5p7/kDWNyJutuQ9y891seRX6eQixnovbzLOL/C0iY9+iP
8C+Rk6h4huLrZ5KiP99rQ72sLb2T6oucYMolGtnvlqkvdBAHqfSek0xHZwp9tRbACoFC1iZh0JcM
ItbryCExrsy0R4G3rJKbqzFTEwEC1zg657r/K+4I7xqwIwN3BqJpLHO/4NQAkVhxEQmiRIeRDK1w
REwZfvgP6vvcVuoKaWcRn32Z/VGvMp2oW4SYLMB/G9Rfxm92gGd88oLucmp4bQo53LY/l93abg3s
zTZ8XL6b4QnpPOwlHnmg3TUn12jSy40Rbc8EAzuorlTH+oh001ABYU8YQABhN48j+/4TxBMwMxRg
tKh5QjOp74PgcJiJpoY4UT7s/HRkCEtSd7N28hckQU22DaYZOultvUTEKlB5IXGF0BF9KkfSr5PR
/3JTN+pDwRW1HCOQqIZFZHsXFPRfARR53FLIEvteoLjWmGlsuVLBhsByFA4dUrgtU28AmzV3t0vc
SQqGu89w1fg2egtqTXjgfFpDgS9ou1Bp0BGrURDYMSELXrebG2tKPgGqyxx8tD+jlDe2J0bBLKuK
EjIqbh82E2l3SsVgakHDzuO4K60e1Cw+c0ZdrpKOf1sRXdk/geREl/OibPauyBLL8pvxrZDIk6r5
LvU3Q3n/mmhp1eChsZB51MLoQU9WYTfWG8CnwJViBmvuN4xpEa/3YzXGfEg2+lD9dEWpR/O4bWHR
KWRrduMvaSzymA/e1DdrT0un+KHQ+ZDLBCjRjp2fzjDzZg9ZWHFvYUYTT5g+aoMf/pS8XCKDEnwh
L2cqWjjuAxjE/fs5tcnL7kjPCRZqo5TxVOTqhSMi0zDf3KvW/bw3GVR+4jgdbbeUjUalZWOJ7K3G
Agx4ZBkO0FUr1/80Ppdcg1GFfsHqN7Bz26Qp9BuEpouR8qVJtJicllahrX+xMnrrH8mZa+tUtV6C
+fseZ1JAfC81M0KQGtBa2YTkImeXgFKkaN0RqDLeNCOW2/ymre112jCqFxGVpFQFR+euJRn767Q6
Vtme7CJUO1XjC9r10Atl91W336HYTTMiHeo//HwRWaupuEMlQ9Mzy+usLKxxb3rFMFRa9bM6NSeE
+qD4fUOlGhK6Wxfvp94aXpwyhZbOHyXmvBETEgQ3bfgqhBYkSsBvI1gjTNM2alB24g8MjbmpBh+Y
GNxACWXw+t0Fropzc5ESWbw6E6nBBBCLf4vIiqZI2zNvfRwp4mh98n5bwodnt16mtTTJ4Re5qEwr
A4Fjx1cpbqCZigiGYt0tEMgS/+mju0CMih9Jj3ZrXkbiksrM4rbIDgukIkEch7eU9K7dWc61W/S6
FB2kNKIftKM+5UH/F9uciFEhZJ6Sj7ecsGS0AuU4HXhwwbYlE3TJ5CPeuqfzOv+rG5plACPd1x6V
JcqkoZWkUEba95UuuLOk8yce5YxRDkMLSxU4CHjpzP5fttMfVwJcmy1TRQCf0cCKKZWEAZdk5pq5
kfsXVKKxUBeQ6gfzg0bc8eQ4LAJEVIQBswoXHpxaCj3jOavYkFP74n8ptQZ31NNnsxuFMEJeMUHH
ZEajArerhsch09UST8fu6xEOO8gqOVtnEEWRegT39h0ZVhQ4xAHx4X7+dv8PrTHgryVHKwbdnj3h
WwQJH3CbQ5gduI4XVSFEaMX7XAq9m36MBArZANsf9cxN/ZkKUcDRdzTd43hrv5eRI5gCub10KQW/
uB57eAXQQRKjDoUt+0RcRy7DAEoH9ubloPLbb95UMAYmePi88TRebZ1+0bRyXU5vBsNziHoyQ/ha
/Mtrbb1OdC7Wf5ucfBAb7+dW1RdWVXY4DN/9DvHLNlEXCy6a5IE53g6HouG9NV67OLNmkcRnLKgR
bA810eiFYkPxHPsQPJQuvPU/4fLj2udaGGcUzs53ZyJfB9Zw4HoltZsoVYJ8yPexAmBz75fewxYi
k9DzQWO1hVvFAdSYIoW5HEp034NgCQ4ym4jbJERn1ohrOlGjVhUla32tharI4L5VFgBgbyG4yJEI
NZ+1H8OWIQA1VERl124NB81vEZvycqx4AwjUUqxcJecp/uONCdDP1eFo6pqSTbX5eS+InSzBGm7C
mH+lWDJU99zsdzoZgaLPDur6KGjcdAmFO4erh/Pfh164njCtM+5f0pqRPmyy0TfFyYswFLLqUvV5
eBDkcoTaFoHc+fXOKfH0uLQbVQDYkngOSuxmJ4xgiJv7eoDysK0oFaaaMVeIDRJNZ+dDGdtERk9z
cFVwINBQ8mr2wejdvoqutG3zNdwFFeOlUG2EUaTutMnZHJdZgsJ+lIer0cs8k0H02veIVEVb7UsQ
n3/3qI0aHQnn/lUOie2r3MZ0yMz+l/YbxFOvKyHPLlw8BSyoG6eYPASxF2HFeHuWhBlP2v2I7hp9
6O9bQGtD3V8lGB60yKQICaw10IT8agCwfleyCgvIe2ssl8gwwpqt4/bumweNICQks9eAnOoGHpoj
yxOqaCqOSV/ZDSy/5TflXOojc0NcRtArbfb4jPngR1j0M/W206m15HelBFqVuD8al4rK+nlJJesg
nlZDoiLQj0NBsu1kqTVpyweDSGfE1y4nelWXnBmoWMXS79B7HW/AmTIMF1FGBKnBPWBI9DjqnuTa
bQ+n2XNVrY2EEzwBJsUnYkCK+0ftW0VrefnCa6oRjNi379qV8NbPO+48laSQ6jBTPzOgCsPKwPdj
lHcVAJZ3t23vP3J6B7+iSt/aZBtmDqPmGgspABZqlI6pfQtM8Sfc9lGuv9nlJwujZwCP8LFMYV6I
Yr4cTkfHw/cGYr0vrGv0qZccE3XC1ITrpG/wduY8S/12h5xn3C5YllqH/URbGVHjl6L4JdSLRdLo
mRAsoS8RHLqNAm38aRQq4wPJ+VyKeA9rAh7OiXREZWuWbEMOXlgeTZ5ux8IHsYVlfyGjVgQIhuCq
HvJFY4SR4lLc9tfhvo6/1e4gCzYjOgDJfJO33x/8/VmuLakv+Gj2KIZDEo9zcoL5P+J06OMxyGsG
Ot52xDvNoV/nvhdSFycD723T7geaPQwUbxeU7DLecx/bc8+CsburP1QQFxjVIB/dzjjR1hNY4lpL
7sDwHV5rwKcdrxDWF66GR5Dv0q8Sb6T901vlpFTkpt6oXuIMamX/Jqber/YvkujdJ6/w6UQg2lMa
AAIuPbnkdDkVHRRIfDN3B5atImbk4s7LaPR2aIsvsEausvdenXfZpd8yDhZCiDq7o7ut9xrcMBrx
IhyA/HBBiFzj5ZSojvqzABCPfCqpfGIiAA1wkwm3Xr5G6/0VmInV1PtYzdoENL51mTQuSx6OAHCT
IfFIrrAGYX/otVdjexpAhueg9mRHo32dakj8F+dh6EDpMbMGyyiC1IL8NNYjYn0blvJkXktuK+MQ
S6XIhJUEVRo9HC/SrlCaTZDa12b0Vvv3GSFHSaqUKhpanMFdGYhAeHjsjlUQOB+3OH2XM2Z2cALq
lWVugcLYTpGsmdjt+XXiLLFw0K3bxLIKSIROCWPZyCzXBon0jAv7EBLN5smHADolXvHQBKff33ld
oqyyuZuH7yKRlxhlzAAtc1ZHMddZFpvq7qNRPLcnXOxE18VrJfNff//WqXmMEm1iTNQ+xTHwc1JO
uMdAM6Ace7712BtqnUAdnBNW4s5CC3wQDd4yGHcxBqDn7z7rU04rnSq8kH12YVvzmBkVeT/rkKZy
KdvhGr5st9AYVbMu4lRZ2Ipa+RTA3EgxVSzTnOx45BcUUuXhyZOFHlkRHcviThydVhLYrYvqWYLQ
4T5HniV9x97TX7Nu3t8ty6lVlIY4uK02znBQiXKQSEOAe1RZdTDsNbeluRDcSpkkfGejTeirS3B2
JJi4a4dyrY/rSYzuywiil2G6taRoiEKy+jYsH9jdAfY2Wq/okGhaefuylHcqwBmXwTW4xqvcN1FE
tV8uVJUduvJDD+fLD57sjxxmOtZZDRS1S6HcfwWaOsJ4ZmTZfRoJW96oR9SjrHZ8dgD2JUk5DpEO
4mrbXdxLH8dJ8LP2tFvFJQtv8ZxqeSfOfGRUrvLGulkuG10sRBacVMSu6WyDFfNs6vWU5qdSioKr
civQdCvdT2Mx2hmlLF9p3GyDJJs+VtEPXRNkyTBhyNYrrLibpiSscGj8UyjYQ5Ld/JEsal1o1jVu
7braHC5ASJXUA8C+OEoI0SNOi1qaWewPSCujCbaMSAo6gvpEY/BEI8vtLV9GL8LjjUvI5JorNlrQ
9ulh4t+AhjUoq+0U72bUevMP7Tf8L24MU2tVPMiZeiDZ/TCfNAijrdx4NpHINLBLS5KxXoc0dUEJ
Ra5UUuryNr7NcOP6NWkhePA3EClQPsgHN9KuLlU/uOmqLlRXyA6xgmmhxNS9vVZOPuG4oO/Gaqjm
eluiQFDLJTZKDd2xptw4UylSxtbKmtgXxd8uRjfEq4GYm1J0ruNJoKOR20R/D4Cu4f42mbw6EETJ
yAejKoI3537p4d5nT2IhjCTDW/BzRk6AoQjDyzqTRyz6WZ7pVT/SQ7Re9sH1Qmqh9FlYAo7wD9ux
DrBlrAC/qvMXOyWbgHQeDZw6rSltCtMTuTjnh14RtxoOS2/Wk1C0KLucvmnKL+b0y0aB1GbOmYrb
kIH2G3zd8j4C87vnV1lsQKEy91ggvdgqvtB0J+zM3Dq91hZObsGbvIR3H5jBuqHyjmjNO0uCVtDI
V5r/fH1erW5NNluxTWfQe48buJKT8cHvIJkB74UBa/xtqzghoEVzsVymLIEvn7NAbGSsIQJQwNKw
DdWqaKBcWNcRw2dO+bGE8ddI6rb5fl3mb6Y3myrdhUX2VuHfmU437EDSrdfPPfrs1DIHojciExj9
RPESY8m1Zz6yzCOlTsRiM8gqkuZ9rc318pRpk6h0OeSXTCxDxDTOrqSF45Plv2g911qgXOPm6Dov
ZNF6WCYyQ1mnFTSKPkxLbBMOG+Kn0cgqs5z2epC+6ZnuzLkodQ0SJt4yXltOJ1CURG17UtM0Uzay
dx4j/jB9Uo51daiVOW6hOgmevbyjO/Zw07xbFGmt1Nn+P0mU33uuwTb4v8qitEPJgUsxxt5DGy6w
NARyG+dV0Yv4/SXYF2KttlYSNwX1E3jaj7tGwPOGjteaK1rjrPbhJ/oas571mD3SLofPUKUnh7tZ
pkYCgqRiXc4kSVlLo6rjNYFbHEYLwW5ARSKcy6C1W/j1vZ0jchMzw5DGGcDuUUGZ/qhrafc+EKfL
xU3vV9Wsab4yKx7P5HciDikRPYmoTJyM85SNLggkGhjLORZifrEDA//PVcBvFKibyuvQVRI/RXaJ
wAUUN8+k980dos0paD1O+8MnLKKBvFCh3i4qv3rHRZXnchCJyDidsRH+b4MUJqBjQM/ApuKN973d
ctrR2Ld9UPFchMsWOOFXGOhqNOPNaXPiRmdR68C65UqNlGNifrOhfLcbCHYm/rlKH5T1O2/hczka
MsV+4Rof29WqQi/ZmjfCdZ8GZ123BsZy6Rwjh7t0uZtEmCCZlxqjUpFPYsaaOGXHycpqqqSyWlPc
uCaGuo1UplS8FEaOZ5pvR+bMsRzl9GooF4p/tL+5CNQ7fanzql33WkQ0Bl/vAzwhDVuu9PW2HBdx
pi2FwnjOqHo0Dic/RMO161fvESzcDV3VkVMZhIC8ZbRDCgjjB/YV4EDKkpOsoQMXCYcw3N91e464
/MLb2ba/JtaK/uWvr9w4a1LV2KAmzxuDFfFT8ZW9Fh8h5hWTEqCvVJ+cKVwH5hEij9ICLJ+BosuJ
Sf2/V3Ig7ww2zLPBPYIE9iEcVyaxGD6jwfbkKsEuYlRi2l6879XtRq5jwnl67RLJ3CAlXt4PcB6a
u0C/vLHumnVdWawKVxydXU2cr34mr8DqOu+ibxvRqTpRT/7XdmLRa9XYhrq6W//DoEucOai0Pe95
CjPrKGI70/wA6g2NSTlfLBRXDyHrGYt/JCyQNH7x5eO6PAYSV0o8zxz5VDJ2vKmbs4CM4ZUHyR+F
2efkz17KSikoKIwM01PN+CkafnU0xfBASdxJppPwGWOSpJw9mJknrYbWTIjCKIjkoApEtIZJIBFR
htASNMzGFVqry3lCI8g+LSS0Wg5jAe4xJadRoJGFRakFN4dcX8P31Lq6Ijc4x/p10/+nJbuR5jZi
NkYuo2Brm0jFO869chRmhys+LlTO+jDphA70M2kH/Pr4IweojpORzZCpVPb8bpB9+7tUYz6+IECp
FVImu8f5USLjcfqb83hx8rVIXqHy/Z/5uPeZstXtx2jQkgwD5Gpp0yQcO76ZInIu1WAcNRZz4JtS
4e6xIqJECjl+izcvz4hlO9reksmlkVau269qdEYNWcQkYLyTWGa85FQ4TT66tkwqlpsSTQQ6TZp0
ilBTIMIynQ+wsDBKTRpeUENsHXjUTBm7VCnhtbgs4XwHViRnl4OlY/OqnC51odBzSKXcMuxqY8Jy
EQFmRH4CP8ZEcHG58OTdO6pFiI84gno66h3JMJdYt7VdKvR3MCMd7wXVqSF+fKSQApbH4SpQCY0M
L+Nv+plHqpzi+aN/61MVEccsoUdvPUyd+c6DD0So0zu963uZGs6hGFGxA08umGbNDIoIq6y9oxTV
PIpIlNI/YHaBDrVo1t3Ua2C4T3EZwdTuZFLUiaVno7j3Z+5Z0MaugWgbpnxn1k05E8VSHoG0e7nB
6+kQLhWKMre0QUWvj/dnZpmy99RtHbGwOe+bTSyREImffp1v+O0swuaDzCUmxO+0vp0SqAsaez0m
tBTaaQW+ykFO0SbJG9UkY0f6rFHOi6+0q5E6n9QDOLtp5kwuESd2xiCuWq/Gy192n53r7SWbTrWI
rM1El6HppEN/tRrnTXuRCuIarkFdMbZcFiJSfjaCTlxOk/kWeobNiALcOQSqEhKsuyMsR9yY5ODc
E0oqXUxKD14Oe3y43OAt1YNYhcIsPZ5P9ntdOz4ImhvVKUEf/+dRM+ctDQQeyrhGJKQ4pDWkXrsO
qYZLOyYTifKzzWYjinVTpoasenahU3deelOjUikEuWNZkHWQI6rty38cGtsxso5zz2UZRwrWISz1
vdcyZYx9OJdOz/pNEit5NdCOxDlKfuxCjSq6RdTbaR2p7oU2tovwylbZoxIke6+Wtt8CTSz9lYOT
v237sdUR1N2DoEzd5/F3+mSJLPiA83fuqk+AGjBfTf4CrYtSggMsRjP2txizCrWVH7gHsK0Eh8Yu
fzHD97KG5GI+nJ7BDjkand8Wbj7u4wBFz2r6cb3qxbl6v66LF+xwmKEK8k6BfeX2rZM/yDp924vP
fbqxPl+pp3OvJw1KSIkOppyQnVEMwsk3keXTSDH7N7xqvSInYsFMKvZL/q+YFuLSLGSvVbICDGPi
jVD9t9vSnUQgvddOOtLPfbttsWG8eSSmDe8A1TOkDsytkWO82n4lP0NtEabXAVUZ4fX1Fmrs3kov
POxn8d39eGqpdYPAgneIBfgUzPdscWpFCc5nDYcvePZJZK76oQBNvMOFlbMKcgWEQBGc6VjTvTqE
S2QfRjNmb9oT8hM7I6xoisQvwWb+1PV/+qgNX+Lna+eBON2W1gCqHhp931rk92Ka1b7Rdxb4CqNd
vnMs1nCQv/pzZNaDTO6dSWOrHdl4SeGPuIy5xKXZfTiZhGhFvNbnGompmmkCrgDkjmojx9bJkfLl
WiR0sLjHq8rxkdL07lLm1q1nTzvytnKF9nOQCvkzfZ49m5uUlLO0ysLo7RoICyGvDYBLVq3ACSrG
pliiTUh0cgzYztJlVsZPDsuvMLIJ9O5VBOrCBt+7OXn9ZHaTNaGIgIr5T84hCIa4XMguA822FaZ9
R5fJPFjkl2MYHajNjunjaJe/WzXmwTgHsv3EzvBRqwD5n66wStYoYo/Zw6Hl+hmkFe5qwM9eTMuY
aCbr/GTaLiR7Vqja+D3pOIaQe1RQ4B+NisL3TERodOMLknsMUSYEmyKX7fbZYCtYcZmsDovBurYq
MMlZZnTInGVzB4KWGi8b39jgTZTbdrHr0CZ2OIzfZ8HmUeyIiWpRMwLlm96lnKSNd3mpO/qxSHaa
vY7IjgwYKDSUnMOQwCepHC2GkPTZ22gDugI6r9FxvNu79cA5to8PKtqAkhYcLzJWAsArCJCnGcSh
+ox2524v7S9POKtfrzCDkJQI+Xy5/9k8gfGHIEfrXetgsEIj5CI3rjXA0UBZFhlpvPHQDEU9+Y92
bbZG+dDgoLRaLKTM8ABAj3orWUhNJEyohjcQj2zmQquk8AeRghraJXfttgaI21dGoFZq2aXytNls
WCHeH/4Y1V/lLxIlKvkBAB3iefsL6dtSBWTvzw6hW8I3DQRd9nFfWUiSGckU+W7TFPD4KTw4B4cH
MSAUr//HvXc36BG54EGqbZ9PM4aXwg/+9rBeVDyMAdMN7EBpoZDxKoR0AIsY4J2T/rvBsJMF85TH
RQ3HzKV+MjfguCGkypTabaOpM1Dy4B5FP3ijYr7Pkgpo+wVLjn6JzmTRw3ch/Jauo67hHqr28YZU
Wx6H4O/c1O9gYhAx2/6BO2Fr4GdJ9+mdsrPVe+I5OCzbDJSnKmpXCSwCEYD+TNBGuKFU3STn84Q1
ypgKvpLvCiIJzNuIMHUEJrUutUnkQld8TzIASR41iJWT6kokOmMFUveRDWcNIBKOijHA19ST4dkf
p0WonEdvfYNHYE4NfopfHDEMG7fjy61LLM/QUvjdSDGXwYedpY4wfxwhjE+BLzVEASDRE7V4+pk2
LNfCVphvH8hicON4QaZvhvwCl8/EyKlWsTHO8yb4wNH0LOmozcwwZwYxVQqotyAoOB8XpUrZnmEo
F3I7XvwwJoTtMkcqHoo+XRv/ypRXgsLSgv9eW1h5s1STUI7sX7TZ0csedxDq/XXM0NcbhNFanbYQ
WaNicOkOhFKF5dQZxVYas02Uzw0wEhC7sT8IKwsHxEhNzx26aT5xHv5dOT8YaSy9ol8L8JzKVMrN
e8K/TVhen9YZK+qCSwbOn8I6gS4IhijzcVXwd4koj6ZxTPRtAHz3ZL1rCZHOc51rX4jDBxihg7AY
KktMIpz97dZZKJQ9LNVMIKrGgQOOoLTyiN2EcjZFoUe22SkbmjXW+4RrNouFaZ1h2c/QOB6lJbKC
W6lAzNVnGytUaF3EI8QbsR68Wx3x5b0mWSDChT3kZ4gOru5R/3ViLlPrzFH0KbrJJHbjLHEG1zAp
EfTwVN2AVEEtvTrMZdbwWpB2odTztKh1w0wiiE+yZ5OBr9ouUROxlSP+tpZLKsbWciS2j4P+XYe8
mzbTONtOLKsSzZmDiET+WELotCqQfPub3y0jYQQNxxKwFK7p1y34sLKGSHzMOSwNDrzKGcqMoTsp
4rFAF/jpO0VsJ1vcGs7V5XSvAi/0W5wpoBgznNLvzFMKGa26DkLCsuUCzQ1rXwqcBewl1rEs8i3C
yO5PGuxyS0D7CbJMz105CMwT92PBeDfjXdK6M+/U/4qZHgT6hK9exs0WULyzy2LQuc4+gNDcAOF+
zf+tH9zu+H8LvD7yqzuGo4FgGbJ5cbwtozRFssq60uEtxzKCTHu6gov4ENNjE5P7cWKOLsDrFWqI
6h3C936yyZ9002UxjTLvkz3J7VjSdnDIGxOQtLK0Qr8ybcB9f9vujMrjdqmBQxhwnEX8L/kG5iNF
+vhNXho4Odeu3yXXQCZbo4jvb8W8LCkKAP9hjZAmPucb1mQhYef5dV7F3FyzJQe2Ldo1qWiNgtVK
QqSZxfw8tgkwWLiyZkv2bUo5ZOh/N2UTKmrmsXxQdOkManxekwOjbx47kR2OEX3xMqRCs+E5QVGP
NP1CMHBRreHSWePcda3RnDACpcVcMcHrPhgWk4x84kIVKIcUi4nHWSkn/Bj/ZXKnL9nIxecz78ig
4Aq0Ex4SOJ/nU7AgdAWoi5kMJXjqqBbp1DbQuT79VHGoCtMXE6O/DInVnUPL97Wk29yaxF8a6A7u
KRvnE0CsEwPB1wSsWzL3LT/d21vqONKJ53frICXCJ58zI7b8NUsVRq+z5eA3xDQxfUW26Shds0r7
tsJBzRc37Xrzax4qAK9QOneCG5sNQk23WRdlsxLVYeFVCh9l0SkK9cU//aXF/s4wgiMJljSNOg3F
4q4EJMgNinENvsqiyjJYO7Wgn2fG18lDXdhEsT5O3X6NYUcqX8GO/9s125Z6O72AWaot8q7NpMEq
vXI3xDKY6oTgR47I/FGwGNcchTrnMka2Q6DGfpzR/1f+pxhw/KSxWHRy0WakT+Gk18aVTxob7ONz
4Aierz41okIPQd88Fy/RZru0KsdC4KfhL+pnxm0sHywceW8gVZI8TyYu+suj2lpi+FbG9nEtOB/E
dnm22FeRHzF5BHXsychUL1lntQOR/S59p4NaQ9xksWTQ8Fa+vtcIf1PCIyMqT7l/+Zln0haJYi8b
R8q3PniM4xa9XIA2fDhmMMJkreZScWPi5NVXG9lkNCYHmCt6vmJsADCw+ZWzBfZS2fpRstHYioMq
MvTzbbrgZxlGQQLPNO5rcpEpdkI6farlJ6Nwq+Z4vy4sqbhEqrA9EndVh1IhBu8gYzI+hweuZVWh
Ziyzy2JtPtIdHpRr7Ot3iHEh/wPd3pRyRRfNDsqBdu4LJhxGEBBGLZodnOdZ6J17beU5BR5tbTsv
sm5Ud9WJTmOigl4pauRxvkTvbcMSrKmrHGK0RDwu0/LJwAoG+qGvz8+5XvNXnl6CJTvW2JEtkMbB
xI2D77Vu8OZNDsISTky5yatyrmLn90/h4+aNTbcEhyUdCA4DWLMTTkkDBlGEJjRv7RGH4bKa4SSV
fMLgpT9lIerLBdB/deLVYH2tN89/o+WU/fqm95ybSsQEJTgCReFLNRDQ8FEEL6m4AnPqGipD8TqH
0ZO06jGDu/gv9/xX3PB7y2/z4LClUPVpvta68jWBs8Yc3B76zytLl2Oocjs9EJj9Wt5B3zkHgc4Z
ISUkNx7VL/XhF9jgoPojybUTtdCY26+AMEO69UzkQW5b4FRucv4jnbuBiJ7jYewaT96LfAj4YoAX
zhdXshO8qi9yFr1ephS3kfPDkkvL88J2ns94HXpUZsbq9Vn2xBW8aYjXEHQwnwNxXYj+DYXF2utJ
jRh7lLNqxe6ttN50LIMpkMUTwNjr9KIvfg4GA58q5ifZlV4BhIOSOIcA8ooufG2fnRTsqWi/9Nx/
xL+yZ1b96CR9T6JxdazI+pP7ChjtuRNxwp1RstpxbjnPZd7NQ9gYxu1maX9mZROYPsFhJcDda2vA
UbH8NBPWmvKea4aciEXY4R9Z+4P7388w1Q0eoZSQXvbQxDiRVu2gykLG4ItfX0t25vocqcqjy2bE
wdBSJ+grdlsR3LH3MYlk1R2fPTj9HKXNEdQCae6LvhRtV1qYhhjqgLl2O+syHLgUs24EAIyYUNZG
iV03+1iJhNyuhFvvw4o28o/3bH60mKhqZ8uP6OccdcrBdQPeQcrvbDITa9YbxAwtll0fl483rUVw
QURwBSrQKGUj64Vb/GNTxpi092MI8Nd5lS58lV2gBcKwR8TcBUfcWySzpBqhz4u7YPzs6A2pNQnn
nZz1FQIbyNrcvDC/uv7bDPFo/gg5hDNPcSVrd/+YT4JVObzjepbofQ9lIkPdtYdm5jJyFL3/aqi2
qJu/VHXTHcCibSBpy7/ornkrdOsjL4KcawoqJosg+HBo85YalBIY1BGK8zvH0j3Hutf9IwOJuLnh
iGkLTFLz44xUYuqzAf6ngrbNj8Ktg+R5zlKguK9oZDLVMWvO2alj/r7lEhwhlU8kazZh3alOZu9m
JTQ6xn//jWq9lFcdvxeT3ttsEff5zA+DucZBIDpQdYPuP42imshufJKJjiWux2KqY9G0gN+pLFJx
styvTxH1Fbaczel1KhA6jx1EmocC7r0cNQosIQXi5KB/V5x0cKsRaZ+NrvRlF3mS44R+4w+2/riz
jgrSZXowU83IeHHJXgl2EY99vGfN/2FZQ8lvfEQdh9fRLmc2/CLOKteRmDOhPJojam6ynl2PXByD
sj0KmrQCf5ZVEA45pZBlTEAiIBg9JVoxlUMrFak+PIgArelXWT2Jf80jJK8yUs7THqf3QwgCfNxZ
p37SnlAFHoAPf0LB9Td/ive96GAT1Ph3nydAsURj5nriB+SVayeZFfSduXisKXgeoZB96VHdWv5U
BGyXWRGsshGDreg6eqFuWi0jgBmnUlrAOXVFP7p66J3KHiirfLT61z96H/AAtX4WI2hHgAE/3mzA
wknczc9HiVvuov/r1SPxq8GuUbRmRVKNbpc+q5odMaX4LjFq0CZIZDHHnX3wvRPbz235S03gwonn
VSEUXd3v8kKiypjkSt37pZkqhd3ryBc7VDUgGWCvENRtBowlpoo9zFVE2MJP9+UknuuD+EsCCM9G
Oie5v+Rj356iz3EHfxsPMz2RErvTxYCIJYVBNa3CBgA8tvUjwCPhNWsO2J45KycRDDD3ugd3yM1v
NJgf7buXgTcsQFc1KAJN55Vw2QNy0t1PaTditIFi90WsBLDhhYE4kCt8V70UG3AEFpjFKOxBPbKH
Pzzgdb49XzlhkZjFotQinCkWhAVLJtjqBhLLIgaCvJQwmehXmFBFdIVGrM9lIDyR+vyBuTZGjNu6
utVChm2+WuEeRIA5tp+TOy1NfYF69HyhUq5FJwcFni0P6jLMZT/SvoHw2DX1Pe8P3OA3M/Ox2fyN
d75tKhfvP/qBbxH6sAmtv+pEqt+TAbZSyFekZBVs5UZdn6FrGkCa3/uu2ba5GD6Pr6DXfkOriOI7
pfxVHJq3ZutwJLLSwHTZ1ZXuCh9iCE+5lApyp4c5jXmm7h6d/rf2eZw0BXXReBCDqO8L6fB7rOQI
nDr3DrmFF0TMLykicdt0gPfiNoolY3ym3QhTyeOVADUR18aWK1YZ5Ug4IgaL4juOQFWpPjqIhAln
dUlre1/PEjYTT++TaT2E7WXSMtcCifnVwdc25tYEhg3e9pF88F8Epa6DOHxljYfbaWEOK55SQnja
1wTyberw2aOSkRs80hptGWlNVHOrKtgzjJnUa1wZ1BhGk7/Nu/8lpH+vFIFv1+F+3w1Wy8IZHcAg
uCgYGz4LG7GiOY+WTSPYlC+izDf/ezUeWjAIv8txBqoCT1rEe1FBRgHnAyX8nDPNP1wTs9F00Xfn
Cxa1EQv4rex5fCG6BB+7gAlAHtdNu02y1VdnwP+BaFqsxqZUYOBDpTrjiIqNOiLpqZpbia6+pgC9
sXox0f+iftQF9/cKcvZE68QSeTRc71DkwNwjdP40TY7Z+BqRy+AZxOu/RpTCEJXYx079vMo1KZ13
N6UPvxt3UkQYDge8kouKl8TFB+DJhDtHL1MVI/KXCOccUSTVC1qjtzGIZZoAAAHa1PO0xEfJByVM
AuOH1qX+l6hHxzczJyNpcUiFgS2kZhz/+L4/w+kiBI4Muy9SzLZOCJvSpjZk09QyaZ2kn+TpkGH7
XyZvoYb/skFYnNWkQJ0xTn16Qpz1cAMnrBHaqyy1l8epxFt9Im8uVNYrRj6JZX++C+KcNNu2eJh3
UWP2XjidPa5VQHqReVK1TMd55mxq2XzXIIaJUkCsvgQ0lRHu/9KeNuKw/A32k27nRzk1UxjPAu19
wRwZBb9yiYZntBz5f54UXDrbg1lJbSCFiILEId1QEo/sK8oji4L/JLlZt5k8BIvA0Blzyo3HcvoO
le0AYlH4q37uAY7thfjmpuwqP19KCqxWrJl9b7TWcz11cuWo3HnN4xXD/ukVbpj6sgdQ3dxZtMfJ
IdxkopMvca86Y0oCbIlhVb0QI5lgZgCN93+3vZDXtpBjIiQFFyqeaRULerWCavQMikm443o6XMtS
c9Z6LRfrOiHyVY2PV1l8Gshlf1wAhJhwkiVo5EpmnpTUgAv91rYUdwvtYb9KsjjRZjf60VKDgpk9
TTKI6w0Ti9luRw/HO0EIayIPU3wa3vta4owMa4uN7qgW1tsfxe4e4y3DGuUVKWJyD0yUsttd+pJb
mSV/iR6xHvOriezk3+2IuSoDVUW3sgZEoF8+w93wrORXKK80yoH7v8PN5lrs0g2vUjG5JM7JPDCB
EqiNXOVUZfyX5CdYyug0akqiPibQzl/cYeObaZ3xqaf2WQkgfUXitko0PiWC9hu7ioGzCO/2EdyE
VFbu56bPyKyzbRMxyKUqZcKt/PparVIBeOHBC3VKQG3EC/fDRnHCSmn793P9z/hKaDZxW2Ta17vU
5zn3Wdy7VqGLw5DUDvB5geNCLQrGcKHjqLtVDG4bCmrPoRO+0WEdfMV/KOM2brDUiMOsSGQNUX++
dbulO1lDH+do/h+w714yIsIz3Z9E4N4zR/8Ckurkab19KkkE4Noh0zQFUCRcC81tt8JpspRiLx61
ao5aI662pxMRip5uw1z2cWVJrjtvsn8nR/uJN8GV3Tdz7ON4RgiXVe4ps3JnGI34Rc+DBv2keFXI
55u7+BSQDyHQOOwnJnzTTXm47aCz6UPUFl4vO95sn9yLAhtMnZGZwmTV7CfgRPymu9rrsWu0vS5f
RNL/yfl/Y9izap4chjdzbcqs5uLQ1qy3puqS/u6AUNZ+d3AOfIi+VnB5NcVpJ3mu9uyU1LmMJqbI
003rZPmfchXWN33e/0MPbccFO/EsKjhYL4TQUI9X5iktg9px/fZzciZiIHVq6zo7yYqtNNEsE8QZ
CEZ3jpUeQ7oTCibpQ8k9vWVkGvqigYGamljTaQTku8c3vhGVkYwrI8aFuYGZcenUAQD1bh7BvWhz
S31+PxJz1YO1vN1AMcQG1HRknLc0qZ2tTFZnv2QmZzhisfGaIYx0bNnz3kV/CAk44EKocwiBR/lS
52VrkordK5F4oB5doHcfi38NrtDGLXIMq+bX64shLN6N5Ujc8HiQSBWUNyiG79k1FWh3Okz8QxFV
nsc3rS4EKFyTzufLU3+IW/kNZKJPKl/u/xwHkX3RZdAzFwVHJmVg8fX7CkT0JHvoBLEoRqeYtRic
wSObiY+yp1nTag8hIdULLSYk3vnKbgPI91LhJvL6YQYx+mhG5EeuJn/FGdlq4jHSrG+saeEgTLNf
FC48X9Gt6sHE3lB2i3SHtQktRlvT12Esf6HJ56sEtJGQnehhQnEVvU/VVRhThlJnhwqn2ePA6Nzv
L1avPtPu7hIiruNXg3w9zpzjdyim9xAprpnpdYAcG8k+Axo0Bj8tG1zbIjwzspILiz8fVk3glud7
OWtUbOYcwpt5wvQDRzQDefke52qop/IXXTuhguSStsl92TqHpU+ym/dtqUxDu07Hk3sw2c6UJ3ea
PybpPPVZI51kuTb2WbqOkBrRhaBfW7rVTAK5LajuojNKQSsEXE36vziay46iaYFKhjqM/9wUDP47
PfF/8jcP1i/I0lxOrYBU/Hb5n0cQ7TdUhRwKGEpWxrsoZA34K9wTSP3Rd/ukXTDYnCYRqYSsuu2L
f9jDxkpWbOepomoUgUI85kZ6iHwrRRNdMW+VjPo2dVhRSfdiLVNJlCRwKHi+v+/VS/3B6kOljCcy
VIGeJ0LtRaamgqb6Ryf0XnZqFTbo+xrq/r8HFvmrvBw+pQz27YVSlLtQa5XsNjyBUm5qDu4wX2JI
pGBGkk+WUqS9CgYqx29/rgNmel/OUC9E59yPt6SJb/lz5qCJTxPPWx/hk/WVwx0pKKDqVd8ro70M
RrZi5e29OFn2pejdSSyTWOkIU78WfHH5Xn4svt49D4/1faa9O62wmKatPiM3BcZZpsEZ2TL/tvJo
505kSam9bE1JM4/DP7g9bcXWM8bXUV0vzPNnRpzCH0xn2X4Lg87O/mOh03YvmuHIHUVLVQpimxb0
CDHEh8Ex3/tK8ZuH4Lupmt7+G/JhgyTMMZ73HkPUBQOMpNMLpNLlYnpf1zwi1ErbqesEcK0VjJXe
rUE4YMyGTuoSrl3/bCzRh6SdeUngrFk7wlDf6R6qvhG9iSlthuFAyw27UGZvVjVJaoRLes/tudvo
OD1ktmARibemfYD9VeptnCYWq83vL/3csfX9KPoEH5IjDm6Uj4MlcpV3SmUQZ9OYAeuS5926LGmf
X0zTvZ5FHOocv5FNZoNAbJTrHo8+n6rUR6CP0sOkJGSCQLwBU/cjlHaeR5RzRxpNTnC0ukGyL8g3
zAr9LLDpmozpv7OcDDI75tq5z2ldL5AIF/84qh0gaRXhUQCf/O6wGa7amvzYC9rso980vVkonn5X
ZeFnkZ6YNf9AKkSDFT98wyofEe0MZ3t/BO3m55UhjjS9aG+q4q4abi6W845Ij5tJX06Qg9Vde5GC
auJ4YTi7aFRGJoh5x19KwafOgiU0llU0OL245nBvY4ysxEL/3CrilDz0XN7PwddhnAsK8ObYEwTj
ydngEcjV7Gts9yTixef/pkPqNwNRzPMGEIgVloNNxSHE/03FFm5gBvdChi3bZKNmu3bxQ5GoN8ZQ
ZSjg29nUOfh0zFRLAsPjfkxZDALkLMSKsJcMz9Wrn0onk4r+sen4pfSnAuSXSNx8pcb8A8iAJ740
6A9QjdTxoYh7fcvx3lAaIFYxfZmYxBaXspfXiQcSrUON0WWNpU9LreGrTnMLZ1bBphPuGyH2oB4h
guDoZBHh4VjftWBRBlC/5yavNDNtN3qH1MJ+Yr0V90vZ2SlcGR3YoZGyI61goFw/zse+7ECa6TU1
YFKOPYk+X3+k7ed3r36rUKMpSXg3lbDZFzvTn75uk21IdFTaVD8MHFeVaK3ZDYapNDFyQipbNjA2
L9njDsG3JGisJggSGPk2Y8mkBP703wRmjTer/0j3BYJzNlMycsvxVrVJ2AdIR+L2wEZS8Mg1B3Kw
RWYi7VzUi9yacnSHJt4y/wob06JBw1xyg8IKE983EbB0QbzD4l2A1psPgbDSxYoH8gcWGAYycS9j
NziKA5qp34WyXiLiHPzIp515XDE820tDbAdXC4HPc+z/hvvT6qDrLfGDkfCH3NxRN5QrUQ6jbkZq
zBXghRRXVnvJ4QYJ9T6RKzz1QxLc5l8kbJ2ypGsC4dg9Dc/OW8NdsVo2fovjo3PHos8zgd2U1Jgm
g3I77WsDZA4cRAd52rT99dz2OvDGF05G4oUDttP2cfo4MRIiY1/FuclYxlk6KdJ7E02MOt3R7zo/
svNEJFAIK6EkI8xUubAnECuvDDeJPgFlNM9w6PtH/uPL7XUWRmN0bcSl9K+r4Gt/JtoDwdUmDS+a
wepoCpVVgTZHJ+DPw0F16oB0UQF1TJUvAmMOgUcrBIxgIaGMtI9vhd5OaxtNzk53VCm8rc93Y7vZ
m5y++C0sFHP3hXCdC5G28kO+Ir+9u8e2tuVkVWvTubnB4T+fOsQsD5TCL61dUPwG/BBCBSt6QQrQ
hZMqWMqA/EWjdUwemXFUdrw2gBIdbjflv7KhF2+Idv8wXLz+aW9qYlYuWfflFYyb+byrEIvs0pj7
mdSTsZAh1cIUQ7xaMlcj8wJpil4ibD/sJvv4jF/55ofiZ91SvYJUpgrmXdE+axda1apCqbJG1M1m
yNyHnUJrlQ/LS76ZcvhPU/+c6ljjUAttyfKz7jWKtGBjMwyXBYZkg0KCuF95kYXi4vGeScjX+NOg
3+R8VYZbmA02OmMGsadZ2SEUFW9DjnWgHjDvUbtPVYeZa0qW76LhIKgd9xPJdpdXY/zeGcUJvsVd
zary6PD6S4/4oM3uMxWmgsprVZEUHW9km8r1OKWNPVkNzrg56sTpwpC+SyFlsOAKBv0vUFJAH5C4
rDo8q6rpUzTIoUhZGHpwlr22Kf+3GmJmlQNRXZ7u3tgoa54fmo4VbCVJOfJS0jIXhuWUzY+nmd7l
xSpwiJ/pYY9O2pwFG4szbg0KvEkrgxcR4mVlfRiHDLov2YidbiCwE5Eb6i0njwWpNz6jv8gORUdB
hbroDomVi0FPH3F6uDaTyfywiX27Anv74fveXsMVYHJk37h+pPo7hr5NHuoe8snb4uVlvcdlybHi
xgUOXp157CTFNII0J8J98K5EM9RrbcJ5UzzevlTvK84YotjBJ6qh+BdVixkfzEaMlIKXq+EmPJQO
hz1UbjfR7MSnZuYbW9qsiYkg/V/a/RgJx7mMVEYXuVqWjLDJ0ILgYxL3EU2aftFf68GWZ2oOlwIr
eDM/BtOLNTima1dhWkeg8evAZNFqGV5Swhh4CFzkXbRmwwY+Rj7yDM4ehO4cjJIP9B/jOtTe3K6o
HBnWu3g7U8k1A2xugLE/Nw+mmEmJe/i9U5Z0Et6OkSTR6Yq09oJWW2RQKC7d8e7WcJziVbEByBr1
paiv556Mj+yxnGaGxGWfKJbZtcy2kwygc5+VULcKNqpc9lwo6NPLnTsfsToOoGfDVnfZlCSZde5h
kuHXtN6hOV+VdHNlpz5BBSK1Ng3gngeP/9ciGBJcdrsBpG5iS1kFYhgsrFROShBcYfTQaPUsy+P7
RAa3Dnqy6cgIbM9IGVxJ6KflsaXkZxxM3EgWvE+/zYtGHroSagG2lgkOySVcI0x2X26nUZY1azwT
Pt6vpebBmth1xCCxYOXnUj7BvKX5ssPO7pg4TUaYWxchXEiwCIHFMeiZ/estvB8fJsoEYVvpEOjR
mO3A4W3BhhJZAoq9xbjxdh8ftPMfhI37NOQBh8Op110B7zCmywKbJFGnJkP0rmqjNDAnO3n6pbrc
NYSwwVhdpbzwtJvjJh2Sth0O5lWdP6MZZXEwS52yWDxKGz4v9nWY1DwP06JNGdLmFWlup8wmffPs
0eKKT8rjCF2HZtj5t//W8Izc7H+p4fvM2rGBT/wC1BJcAQkqdomxoGmZ3iV8yQMsWJBB9Ae/S9xZ
2vPCxwqtxCp1To7SeAPFF5W90P28YZx7XN+A7djNb02QBQfe7uZD52Tgy4P2+H8ttENN51xZbQhx
5yrT3bT7YBr54P2I62aX3SHUY1r9BUJD3CasVl1LJaHkcOryoF1NfCUwRVUHsdd7HpFbT47fQxxu
o60LBL3rwn8gdt+xpXkPwI2jGg+LAWCELRYvs3sN7RgGTEBG7gNcsWA1NRL2EnP6xhOUmU50SiqH
Wt/hebLqMTjkdmT9trD/QKvEGG7scyrqslaZztsiLau3TkyyHzWqBDEj4YFbTWokAfSgTmEnWK/L
bMDVr9UXUSCL3FD4kJzODV4JqizB3Mr/5eSokoYTNlwVmVoffRw5hV4s+k3LS4dlDb2tNDG7wd3v
L66xREp4urbtrrPPKYm7tVcJGENNlWrD2jLk9+0HxEE2klyNLlsyIfsJDq7jxJ+WDNA6Yki3GbX3
I+qAMAHnDXZq7rZxgtsr8w1bPSNl+Uzn/4hVukmv8BZLcDiFnhIFDwTl843Atbg4SnBll/ndIW+D
juUcF2Xj8MSB8r3HCCqz720XYfHN5ockSdxD1pZ/pCgYblJPJHclzySJcx4FVnNtrCW9NwUnIsfh
7YcXILas9caVHEqNS7Ois5cb7potDXnGt5nTAulMROkTjk63+KFDRZ6dGJ2JpRykxYIeybjRjt2K
zv6w2KS5wI0AHVKx8rPvfr8qsuzNXRk4x7loSRqOpg6eQ3efGKBF9HX3ms6VVAy03Ndn2nbk/ZBF
DBqWRvSSXNpYKhiHYXowsbVa5x9lmpj7cTuN4wFtuxsWXiMeq7FO3lA907kcDdfL7zbE6KsNpYs2
jTaYiYsS8vqCghlbcfgPz68zByaaPevFC939N/tYLiPlK4tlJKFDjwgqjOzEtFeL7U1rWwn9LctH
qf5uLyy9i8brkYvbFBGU1FVQinXdDhKZmFTHS7Z2cGMmE1AdIyWmrFN3uFs1flAP3vOesWxFYPM1
YGTnY/ffRnbkZx7usk6yfLaDxTnObhNfLeFkDeO7U+t7YqIhTNgFZk9m+o3TgGnhScmmLf64DoVZ
EWwwGXA4ZtxCDTOF8x2GT12UQjISjnjHz4B1FW21AEWvStKcqnpmToE0GwTw8Ccwf1Cgq2d+Qy6P
UBuB6e5PjFEW8ZJaDXXjVhjGnxFhBYPSlQ5nX/YRG0u1GCCG8mB1yp9RdqDTgJeq8cENQQmoklNv
tMUh1cyCdeEhl8IMSHYEbblZ5MS0f2TNC40C11DMbFKuPBoRwG5cHMGt4kSi1gdngARuO5/yA0rF
UcurgXS4dgyHPCHR3/2X7C7FFM5FI5ngIo1iLd3J7MjYe+MTOKb2w0oALifxGVcygxc/J+dhq/P5
cmZATEQ11Sg3b97rFrh95pRu4iVWfLhO/YqsgKJ4GS8kRcTMt/WBJ5j9p/thqR8xedICY4SQmLIs
FoL3fnFAmyG3nzHnGIK8r35jyLcFnULiDvavpoQyspQfRYq3g1Q/T2qljl6RvDLzFJGdU0MEMYNN
KAUQNUlvQKa4EWo2h6G678Z7/eyqR43aJIEM1epOYMNJPtTmfygjPqayp8Dw4ekcrqVxXcP2kTdu
3XACxSrsTQZhAr5LUFZXCkLRk+R0kAfDnjfA/pa9fHpYH0bqjsmZwebcb+AmpUJGn/Or+OG0lVer
32fH1SQ0moz/c1K+jtyPry1LCRSP/R2Zv4g2ulv5ynb4dUNcaXKDNvGugkZ2OXBm9pNRP7YB2n/g
p66Ks+fPUxV1Y+qnPrDwJdr8Oc3ChlDS84rH1xfsw3VxFZwx5ClgBCdCwmyjne/OPX1gyXFGFqw4
f1RTGwI94HpYU5Cu6zh0hy55tbZkEcnacX+6WsfDghbZbXppCF8wk3ZUrMRfYaMjklQTxYtgMef3
PW1Oiq4jDhWAdXh9TjuukKe4R7JDkKJM2P0XbQrxI48lAVddkoL5nlw5V7ml1a2D36j93LHfhP2v
lLJeZwKSWBuUnfLiHBuQVlRWeEsWuMLH3y+HKk8AR/TMapYxb2c2B0dncZwPP3anQoa+6jBB9fpB
KHwwfxQReFmOwlguSr/pxuUMFSyqju5ZQ2LeQ8VJVDfTo4MsfLOd71T6AaYSSFdf/MhPr1Ef1LGI
pC5PjOcvs8ppnGv/FbW7M1WhRqaBDrXd5kRrb5CN0R+oVcWIQUFJOhfinF53RoRYotVKsGbZtYm6
egl3hm0toku7KOjIiuIQ/q0u35hjru+QZmsFVtuS7UEM2nEuVBifpCzkA0GwuQTv7irP7lpYEBd5
bznz20sIDZEXB+i8a9erK5oootjc/BM6lx6Q+LniYqi2j7v7IF1ZDaqMA281KpccDmpJ9TOX7smC
eU9t1pPaEjx3u6Mrbxw7LGrIXzouev9OhgSp8J+jh8g+Ubg35Gs2aE1Vrp3gupRe5xw2h8hr1Tuu
M51BhVmmoJe2LYnixl/ZLVxxuU0funrfGFZYKjTaGzLIquH8QuHtBv6wefiWq/KRkBMUubgQ8Lrg
6kk9rJOjl6Mx2U7NfTyYIRHMpeBu7FgGBTt0QZFjBui5B/HEGoM5UR6TwB7WyCW8PumdRPpNawkM
wuNCsxvtov40YBzYWbmLNpSWPfa9wOKsRJKNNTw8Nf7eS75bGVgggJCoSGW0B/f4oti/fGnlK+zP
1FhtC7ktiHEn51hg8zFajbTdM19+3kiVI7nzZYOyQi/Qg3Q17FhI3+xc75vgh1nE+Un8qWZX49Rl
ep26Qt/1YKAm4M3j8Awo9Ha6BVPT1+igBU3Z2amjSrnVkzdEbtraGGtmWp9ADh9l7/XRs1GU0+kK
nAZYu5c5RM/S3N7CI6uxMp3Rm45g02UBb5BECXH2NFeItpoYsRB5hnUERK9j9hR+J+mwRDNbxy3w
LswbNCVfVFcvd7n3MCw10MX9GMmi468P3bypOOScExmuz2MdZ8RSb+gFmxhhJdaYmIa+Q0jieVZY
JmyV/ag+oyc7hUSQAIGaH4H3EX8VVPCSgVwkapVvdzDlOmsrwosOyasxQypTDKlu32t2kgBOuG7G
TiEJJGmfbtB3YOxypzE1sMZPA6HxLovasOiyZ5S7E26bO1+6R/vHnQ3Sv9xbhHqeDNmz4soaG7pW
BpNGeeYLMjKOJLhgvOyN7391oopKt335/XMMCs9YOeiIcTLXg244hDwMr9dHldYSZBSMD2HoXtAD
hjHk30PVta0gouJEgVm3e1i3IOveVDzrZ1+89elZNU2LipS2zOGgf65KCkD3TbPUNRu+JxwHCA8q
lxhBDmIz0uDzcRKPEzMZRq/SIKpGtepO4yuSJba94aIXvUjKqw9aah3W1A08TjBgkt7n9hBSPZPB
LsEy0SIUHH59AX8vrWfOcfQWSh6HdYGivRxXHUPuBm+DFKyN0UFPorzioIK6brGWZ06ca0iDBxYD
RRfneDUGAqV9KZcT+CuOBPRBYB+BmXe4lSSTVNST9xG2RZMzikJ86tXWw/Q6FkpOJTiMa2wBUS2L
9FTjxOx1SwH8WurdrugVyzYQnP4MFrHUKuYIgbcA1nuMIbtbPFmaVgQ/tzRUUDmMQENfkAxRDLMH
+rV+iwVO7AI+Ox6vyEq9aHUzshVOtNv9qyHSCrIoF/bDc6yIdx5NqpGhVHwEcf/SK492P+/AoBHE
7eTSiAGb7ftSDUMN3Zxv96zFjGGewIKk9tQch73xXNnvEMxaU1/Qq5slE+Y/IQg1oOMf5tu7FciG
9nkj0IlQjnXrXRkggKosBGIPetl8OdBS6wgLO6AHvKaRNR2zeheCatJaoNDWKkMcha52qABcaFIC
9O26uOXvPNe+gkIunYq1R42rcGrW0BAvlLtK9Ubmcj6QlRoLRs1MsbAJ/0M2Nx/18qZsh2/Jy9sq
Yxq9+VXNjTfJCeH+YrLarZFvkIYSLvJIjJlRewpL3N6u2duYzsehI1Ep+xmStu3LHv/49bdKw+L2
QvcpE/+DP1+C324dYoBuQvt5UJR8CxdqbQhAFheDawTGo2vf16w+KmDn5wlg1vUwL7Z4pxnmYA/y
bv8u6RE3yLvOeebAWDa2drayn/aWI8YvA9q7aMvHTsVVDtUE4b63SL/QjVWqPj7ynOL7f5SPBW9D
4qoxuChgCk7wmP6OCgQp21CsYzb83A5mhyh2d5ULN0ut7N7wfKbEfjH41pH8uQiPCPg0bjirKZZM
aAllGWM9bsJKP+uoWrAdne0LUhAaigOMxiN0mfwDQJUbEzfOXII6IekCM2ULRQwRUvAWX0QyxXiL
DfaFFxELbpcZs7im/VFX5akEYKKLE2lA6c2AE6n5X/E7vVS7+JcBpnMoZGCCVUy2BAnhaxM43rEj
tmCK2DG6iM4zjmRNXCG3GjNv9tROIdYuYCZYB28TboKt5HLGAi2Oi7qZG7Za329F5gDmYTd+f/qH
/CHmAGevfZ/XxcLe2mtUyZBNNwGBKg8Mr/LVRwEn6O5Ja3uERNRvjHIVkcRD/jic9+IThC+bRwz4
QeZWOGR0/l+PM8fIPATTbET2lJF2ebcQfmVOxRgHRKoQV1MJgljAPy2YAJfL7+xNzUI4fbIcsbe/
9JDXFdEVsjZG91CfRy7JMQhc40GI+UzZuKaIjkssZMNfZ15mzJWtvbd9ONx3e++epEpL7m2+ASvq
wVB5OjD0oUBmwMaBTV8B89KuYLa+lZCXUD1BLZ14Ia3tmbo7srnGAC4nVR7BQkQL8XauwIQ7OCIw
S2IC9xTHcXfEqwoYBorlLYcHrSiUUb0xwJ/75oJCNhHdznVQhZcOsWizTVjk42LgORduhx2YrTCy
6nZn2AF7mnR4RKbZc6umriX35S+ITesB35UGTfOHvBryxmbHG5/ZeLb1ykCMMID4GlkgqH8P4i4E
iPDqoO0s0jDuSl0Df5RIHlyYJxj/qivgDn7bsRbgt7e33Q/mhE1Y81gO7/MdkdhMsbRaT/OU6lbq
52y5RKmOrxHOrMbju2eYPK7UJWAdUZ2qIHTq+VXcaaOje9d6AbHQCdXbFUFrPg3JkYjd2L6ycc3e
3xUUb4CkH3SxsKAZ5O8mSiPNvz/ZyqQWmGTTF9ErzoNxZBeIQT7mYEbeyu1exZ3xo4eoeXnEjEni
WNuoazMSOBaB84Xo1G4RnMmyqek5wElxxWM3YiOFruC1thR+BqljjR9CRxL+Me3Y2S/DcZPLO6se
Bn5VBhzoKRW6mBDxEStcQbkUVzgQHfulFeGKmEG9JpwcpsX6c60+yMN4x+ZfHN3Fxd0HPNzBt4I6
zZUow2vyaypVIJpn8vdTa4s/lUyu6onuk0+CCIOxWq2fJB4YjSjjJjybwcKT0tor/UDXEpVi3rX4
O0bK793F8Z1sSWDwWKb0SoNY4W6zZbfpmvEDPDlhU3FALUTizUSpznYkzcaZbZr1PyL4PQV9z74m
raTBEOfFdMq7yISfCPxdfePJzBShJY19GAfYF2DqOx5KImq9TPoI70j2WPBeCcnntFGBlMuwudCF
W/X5gGqhgYKBClXSCxTIb/OPPT7AZpYYOsMgwSymGWH9iCNU57ehpyM06czJ7KiZsUpnh/khLFGw
OU9rAStBpVJ9xLdSaN56i8jj86XQH7G5rrxx37wJRIUqI+GSBgppRJHZVMSpL/1ShaMqumD4a4Ln
KOM6mV5saoxvA4Ths8ntQ7MF4VIP7++ccf1VoZIxrX2QRfRRpvJXUT61gcKKJSSPWBvQ6pF3XQDS
jkT8SGyGSscM3abLxNL9xpqI11Q+UGebbcpCCZ25pNUleXNy3Ilm50+s8vo0u23JXHmkVaVrJWnJ
9lGpTVnhNWP7dXS+50VntYI19muva3kzfwisJN7O/W3tQ7YWxe3+WvYjr7jaDdP+41rExkFdvw1s
ZpyHmXFOIwql2EhRXCh0ZO9uZOEbW9F8z69s6DL0aaqYdFn07QP1Q2uHuUD2cs6DUEcrSRhzRqJL
fZgia9f3NUdbXtWXAcIVUxFEn7B7X75kj0MGvjilu5p7n4tskBUI3KPylOIvvmFucKHGf+Q96dJa
GCgpVJIpAq2+tK4foO9DPVHDQ4k3eJ7Q1t2kC2woV6b7Kyz63Ttg2+3LGQJsROKhTs7Eqkv5Tmnp
6Eb2SwVGHcT08IaQ0/W5aDJ6U1JhDOuhwh7UliffBIors++J+ID/Nw0VbwHLT5Vw7Idt9hKmsqfe
8RqZB56rRVtRsKwwttgGS5TEWg48Lg9F8PZMQrraHIghz2pl84GWMz8FcdUY7Fxsbyv7XuWgXtKj
hXqtqecrRjVYr1EqtL96fIsnAI8RbWPnf+9o7HdVtJCCoCLGE3aq/+KfzcgyqCO03Rntj/hxKEQ5
aUXRV0tiNPCc3BAwYL2AB2UPZomZowEmtriVSSInt13SPEv4CPLNJnYfCJ9RFL5q+MiAtbKJBfMc
o8HMm7xGGVkOCFsnu5HGx//h55njrI8+sozPHpDTYU3z4rNeNUGzMBlXa+vQ1THDUpiFDUWE1R4L
GLcQftSfHtI9MQyaJc1NOrqCFaX5lJbPtxIROTFB2NqKCdmYPxaFXNHTBdCiAs4DP1PQ7CIJkHoa
/sk3z/vDji/02lTuAfI+2IJxhCdfg1LqK2BcbxL8+Jk3d26cWiR1GX/NZh2qXq1mwImoWdyktNRw
YlAGQFjOptCoMJ+e5Z2kO9kH8389s1LQQTtW2bt+REbD2sc7QHXw5Ps67SMZLQ7PWG4d6NtNE62K
gu1UP2Y6/UXjwtJbvUr1WkOxOPl50LkEQWUyzqMNJhkWVlMTa5XyOWgdF2a9fMWOdGgU2sHCDBBF
GGLQktWGeIlu/qKu22PEV8Ok/Q/tdrCu8hPz5NvvRJqVQ0YpNfNNu0OIaA08RWLDc+7u+eGqeM6G
Bq2xe3OCjjl0r3i9lVDbyBJYLc0LnG3sL0f+Lvty78MiIesc2A2AUTbk56X+VTb7cLjrmTfKdyCW
Opzh9l1dZbFanjBC31wcQyFdhNuE/w5zJ46uv04UyF2ynCkYK7hVpG84XNp3li15mgEpDrCsfNEN
S6XUD3h09b2/XaR5RQDea+xXGHrCQXotnE0Iyxo8aSFaaNRboJVYHiNNP0Am+A9P3ZqJjBUA7FYi
YcOUh5FvirAaMmqYYQXSUM6KGzkR+3Njae8HT5pQq1Q1lUITKLYzmGl63Or1Kmyf2ybzMNe7xxkE
66wouE67crDLze+chLOKpDG5UhuFfhmvZyHQNwhpc201s2869V+D3KGPpqv7SPnvPYMh4B5ZcrBb
qn6qh3cNVpPHSbs5Vz2YsCLehFL891KFohQ2dp0SJEui+q+YPrYYe/0Ncgfuc36zWMDimv0WuKJS
ib7jn0pEWGPL6nKnwcnNvI3RvjQNFhS2VAaK9+elR3QlFH0E3HN9otX1j4fH2Dfq3wFxIXLp3IZv
bAF+QnxZcpso3vM3fwu70ad8EJZqQgcs/OeSoPeSAFuj/sXM2LuYxBhTdEu/MXtwty+ShBGuu8B6
++asCFqXXVXXIU8oPJVk0ZK7tVh0wR7qfFiD/IYG7Wb9o2Rca7ve4u4Kwj0TXfm89vGaCy380rH+
VBp8RhHKF72gGnwA20M/kfoJYFxQdo62vwWSxFQ5or5idt2al0EoqCwzbdpZCWxRg65eLON5AzOf
PLreMdAwek9HpPM0ZzlF2acP5i+zEwv6U3FrMK4017lf6ugQV5RUqdB9VuGq+RMa2BOKxLzh6QVn
gwx/IA3UEaPqBfYgUrcyhpxGSutfgl94EqjKqP2E+S0NuVoH0WCae4qcpXN5BL1Fn4GwTUmr5cyO
K9wrs91hcDIEbjl/6nXkQOMrvKg38+Rect0JDdPzicZqZRoXpXHta0VN0slvexCFCpEbSSmfOALo
4ieL+3YQ4IZw32hY7aH2GJATtuw/4rUwGmD2cR3kfBASy7Z121iF9+jwglsyeOlu9M8YtMiPH4eu
CW8gQE60gGhh602MPCZwXATVqfEhQ9L6LpBMhvlG7jhjcbgGmz3otMAUw+8ktSCy53oBXLrPq7qf
JZVWBbU0SN76IehLdavPEYKAhnlDERuvqYvi33+vF9PmvTddudg7bDobUHkV237ouvMaNNK1TZtX
17MNW++21ohvZshIz3vrbqwnK7HeHF/PtVOLz/8xhFrjV3YnGg9TGf0RnsbQWtOlj59MCwVrGPMn
MASBGjbp+pYJ56ZadiQvsh/A3YfvJvtfHtNZLX0g3LXknRs4JHlt/ua0l2oGkFBiVpGOeTxTIQpP
wr1+1pw+wEGIE0tPR4UTwJ8zKR+2xNzGW9yVUfkz0/VvRULlibxGp7TKaiZPv8heUb7mHLmZEb45
KWXJp70iujF/CXCt/UF9KNZHbWki70g3IzxKRtcYOY8SNHZpywiXTf4EciKSyHgweKBt9x88xbhf
/x7ZtmwfV/zKul2PXtqpAbREICwSZAhVXOFIlxZWKka7eKGDwNDVoLi5BOgQoGRQZfFdK4IqmUJb
S3G+6HqtzPMTTtL9lXXDdJ46Zl2JTzEhaXRqtY1sxfyYaUfajUILi4U0YD2K9ScD+Ofps2liAFqp
ANrXEvKwfXS787XnyRKGWRXpJxM8RjzolD9nbyhHEOsbEYWnH5OXJFwi60kllEhfhJn2ad2hA603
b8n/fmyWJgkvVblze6KuI947Wldlssn5HJXYd+2Wk9l/iDP3O8HRPq3WjqFpbzrgw791ujoMVc7J
PQ/bL+ycXpCKstS+Zgmk5NAWQm4t5es4W+Ml4tPjFRfaZDnboKrzaRZBaRabOwaqWRCbu8r0YSRt
Lnvw6NUR5jD+qsWOMK3eyNsRy8AOQcY9yVf5XyRG9FS6wpvO0pb3PLmP1JON7XjF88Sj/XIc/nx7
kdvtx4Tt0ugKhLdicnxfQT0hApAcus2sgHlzGY3RC01LYlfvpn9ZJaceKnB4+HvSjAecPmEutgTM
VmCVWYaOo2EtJpBm29+zduWyss8AVslpBU09rQ49V3qIPNxft2obmzDzXE2xtpC4kLpo2ydY9ENa
RRHTOlUpAGUbTenRURvZAeR31BZbNNAwvIZaOasMVwmB4kyhOHzFaACWHBZZnuAyFiMrtWV9GVsS
PbGyMkOurjBJOgUjkv01EtcwDYv9in+Fpq+FsRUxLMs0de/pj8ZQ8jLCvogcmexmQ13Zu7hvd/JI
1hFzvbjdwJ70OjtZQ2mkcoUOypvCppcWFeTDyqLXfaMCKta/VIsJV96wVSuoNZAcaBZmJHlgqOFP
HJje6eyPjjFCptsRRlDX00GTj6sDMqDgl9Pk0BC2TBM+bKOScffwVM2sSJwqIylB8Rxx+sw9aUbv
5ruMtEn5Jju+EO3C/B8ELL8V+QTOzh+cx7wxOm3WydStQF0Ah+P2IZgnUW3SazZ9CCXpNzzmHuaJ
pT1Xd9JnVxaJ+Guw0nJFmZxdyKhBG4REkuF3Wq+k/lSnuCvp4UfWq4CShXfGVHcgQXnH3Zf7LHkd
j+4/rHbpvMGPfrB6rN6FGtaoCSnXDynLakgz2OCh+XaKq3SMnh9rv+UEMbEqU6eYlkWVK6nxQX7Y
VxdAVyaYhUnrEu2KFJlk9lafQSGrtokp0YX/t9dORNPspSgFjypqoTmhgNsfH5G5O1msGgbkWxjG
u1dNN4HzNS4ZobucWMoVg3nno6uchcp4yw68aPsNi6sZZArwXV6kx+klsPur80c8RllJzgqxcy2B
mlHo6jP8GR1UeDtOumxKpBcrp0cEgqRQrQGJD85riFoGZaWHRd2rvaEZuE4QAsjifnkUs2TS5/gZ
FwyLLk0rQZTHtkeHCvSSlgOxTQ0ivp2+g3bDGzXgPswFPsp7n1zDzJdAgts5ySHeP3YwYYZnPyt3
7oH93ibJ8MZDvIyPn9fDStpgMdPD95s/L8zp9ivJxzttF1Q7CoITKMtXBj2lNZv4zBmm9lxMOXCz
sUe8gPzypae8BeJXjeEwyMDRfccHWTXjHBBwPsIkQOo+4bsR2oJgvILassBoy6vmm86Bq0XEv83D
NFkoE3jah+E42Sm+4spvOD3CSGhdZZyXJsnRvmSYsw9FzW3vVPm/Hu+ytHzu1m8uCoZQ/39/71F2
z9sflcLMW0nJg9DkIimGvFqxW+RdAMOWOh7vDDDjVtHaki9bvW2FJBXh8hnBG2hlUUWYVkiwpTOL
GSeEp6UWFZV1n5HvPbjS8XAx/ps0xu3iDx4WB95zwRFm6GjK/Z3Haty/auNYpxSD9eDxUvDVqbaB
hCj+cHiDKfoy3PUXV0TPH/PdcPr/bo6ZadpmW5Xz6diF6gvtmIsq8IcSpn+8MuopCDBFMgZIdfbe
LJ8LAI8PB3DPNmACO51P7LL2xOtSaWN3guxgwNTve0u9x0W9tKdDOCogrF24P8B34jz1OXinDHSA
Afiu30QgurljervaymuWRRlhAQqAHulX3ZzWOnKeYzkm4HaS4Jmxzia/qm+L7mDsHdXZGMC2rdsE
e6pywOJwYe7ct7X+WnRgLwNAo4kb0p9c0FiXnoB1ECvMcLEZp/u8vOot6Adrz1b1Cy3np7txqb/y
abf98zO0XwWHxyGG9DzIzMtQFbW4lYq0QPthc4s9ogJdMZDRFcpCFxzEawX2J9Bg7B44Icyokf0A
ZTkvw95IEYw2Hca/WqKfmVGvmAY8E4PH3HVaVElwg4EK/FsJ7m0JfyO+lwIPqrgdXi4eM5gri3l5
bbIKexRkAkYjiZnGp7VTzS4BEiiG31kqKQv8yJ88VHtg9Cjf/9T24hrkK0XNVjU4SZxHaTtu0K5q
rwAtYB+FII8oW56IVzj/XmRTAPVLulO9rVa3whzRUxIzwgi5qV+uifrtTMgA9A7MM4+JBSnx7UKm
JRbbgF6DciCKF+4SPzvNxR7UYYeBrowCS/9SFYKOXQjMZNXLWwuDEmqgm51vk5ss88gTJVhiszgI
dD94xJYyWSlu6W9X6xMSAE1WWkHihUzcllxawb1CBUN8SUgSUblV6CtwhAKDo/jH2AHal5kSxSaZ
eXtmWjPcqYZi8h+WWkudfGRiukLerFktoztXj4V737ZBN49gQQvtKRdu4XfNNITekRCaKyLpjyV9
0fOuC+4QrO3lFnKTS6Mj2DhmDE6HJXIqNjxS9t8p/EO/IyWR5kkxw0aBPtQhzoKR0dKQ+I0+At4J
4UU/1q4N2X5v+drPBUBZeCqyvG6HiY61clGII7F0FT8qJocOPKrnQ8u8Vs9cR8OrKht4l6PM2dXx
HJPW13NCItd50TEPyUoD10cBgw0rgyYqoUZAu4Gq0Tgl1Ef6MR4flG0599gieZ/hKfw1sXlO8IfO
ZQ8gKRAn6wl2dps3zbhFKnCnGV4sqexKvYheNqepQ+JV0m+xElfCe71YVBDC20N/T8+22SYs4cJZ
2WV+QAL+CV640rZ0eET+7hfM6EYW/bI3+tll3+5P7ku7+Prcu3CNsKor7TEXZ+TXHplRTzDxzHtG
8n55ib0YP22v+x31uzlJqJxWqAd3yP/e5eC3+n1ZBeVeSgB4216ny4ThvoCfNnL0dHoygTiLEttJ
0pexJf13WmCQ/jk1aSt2OX2J/rqLg5G7WLyIUo+ZFPZYiECKadH49KE8u1348VhrIwVpErXMbBxA
U7LsWOovFEVTh6gom/iAklwn6FyYMQdT2K0JXvTRzZhEjJiikgBVVC15Y8XjW76r0q9OwmvpHC7l
X5SHhPO8Gpvt6eA5ItGt+tfLw7t6B8U1Od6iQ9rIEQx+XNNT5BOIAtWUb8UMk7mga9yEZYxnUNo8
nowcoYh7yzYdCTli5joz6fJu0DRSQ4ubdaOtlm1PmT/OYr2DeUBIP/JeoHDtUM2NYGypPfAkZzCR
7mBVpZUI7wKdqfxwjy1w2SV/GKC5BS6t8kY1kG6U91rnM5wejhWyY16/UY9RYxkHVOy9u9xiskCq
5NNA5p8XtEEgnzidQPdn/kdDzmKg+RHxvdQBvscwS2zQAHsuuSgHh0c5U3rPUS2GcfFWHK4elIK8
ZGwZ6wZVbzPC+IqRQxMRT3EXlDsjpw6wwXHIuejDOYi9v5Z5DMWpmqpROaFWKn4M50GArGSjFgDK
uP1U+bF9GwX9oky3LYeFtcoZpmLRks73CEiV/Q5QvT/a8LHXZq9qui2TY+MkrUsMQCCJ6+ddwzq1
zpj/RHAA5RZdg9GI8zB7bOkIaa8WcrZKYC+H44B8jgGVAZDhjXufE+u2m1tT1t/dkCGmUNUlgLNo
gaMimLQ7pae+AEBE/DlKeekqODcDyB08GL0Ugilfb2m22rvu/kvDKdDoxWa6ZoIzHaHLkPb3z3EQ
85Hxgppidf5dIstvEj0C+5LIbWPULyS6pU7p9mgxWpBPcA8unF10EyFTFCwb2R9pyIHVCJmtO0bL
bBC8Yxv8BVZH3g4YJzz2W/QaqyXwvdgzzNV4Y2+HS9MXFHD022N9b0dLkdac2jichJxbrLPSHN0B
EO2jcdxASWAQrykIiGL14Y9d9xSOWs4ILEd4aYBAeAjUqwoRW7WRqirs9EHnWp/zWk26ObEfVnzD
CBwz2ZQ0eKJ63q5dp5ME2aOiuYlAmZNCCyAHIYqrinrTevGdR+e8p3jD2plk8bF9MOPWUuS9+pp6
k6+xkZ0yswquMrOCD16CACPdtrhBO/egae1xupP/kiYEigzeMcP4YSu0YNLkoeOD3yCPunMjfP9s
deEH9EFAPh9psje/fMVkChO8a6XG+oVmkcIdd78lCG3M4TmVtg7K9OGL9n3yrIsulmkWmwlRV7yk
ej5bvCXiqlVbNkpuCT2lNbO5+C7iVkCR2rWuUPhVmhNy9aSjotGe9+WbN7AyEqlNSDSCHfXUGhzh
G2piRWgCT7Y01uiLIQSrX/wyPdGPS0vIYQiqVU0H3cNs6HgNOgxvfrfMzT8RJ1GK4bq71dMFZflv
G56IcAPsslnnFfCz0rkszTlhzfIyi8nsKKcx7A26B27f0ILpg8kjeo5jzKGxXkLr/9n9IclvQ/it
HCFQRBabWrycYkjk4v+kh7KPppcFZo92gP6YFhJTpQV/QS1HyR+q/l+AlcJBrbPJuYLLGOieXY8R
c0Px6W5J8j3/6iDKXiZ5GKP1+0KknkZrFv0cwk5QwOurn37ClDPzGAxfHpequcUt092CiZoZANrR
D47HjxBs+Qbi2JSMKwVtpRKC70HoAahQCK7UWUAp+OcCkujH08xj6Ae2/flxEEZscflbk8kuTxdw
x/80GBBwV8ZJYCN8G9/8Fpj+G2MmFpazaIgv3Xg/g2yaKICaWqEDOejlGCUuwTEBal7Y6mujHpsM
wZ9XDld7D6yWpTGnfqZkj2g56PwdTwnrShG8eS0/2jDkF8ziARQcmkdKIoB5/mgMY7DQBkx55u05
OCyKGQdtTHWt+4UTMJ/pD3vPQnkp4XO147kwBPHREs4zcImWWf+45GWq94JlSPZbePYlkUSKxxOv
M9N1YszLYJ/s8Q04E+e62qFimqVr0bSb8l4GF8c7adlnoYrYCnuOaU+qVRbmLm5LhRLPTaVjNasZ
P6ZnO4RaVNTXLur0/CLLd00CniaawvUI+kvzGh+XLwzLKXqBsVDyM2gejKC+thEQmZNgowDZXUmr
3I+5ww+bXB8ZKn419vNqws2UkFTWG35Hc2fhAoTLLRCB83HoY7wm7TBwMYQhb2TkGniP2Z/NGUB1
LWhre3CgH/Jyf6icnogXYCL0+oZEaFlQJcEQZPjT2g0q3tTri/6RN4Uq8rg1r3Z+jlqe1znDuuRu
LBK+pexfNV5kKPWb+5G83j7K8dyvs4F4h6N7exXUkmLHliZxVGHLjdm3E/q+SCGhKcJozgDzPmvY
EgYvBP4/nIVeZVPuG0MU/Z1t0jPjcOfzegDDLWOOMOs0dUDa7pOwOp3jQiwNfF11LisMFXaGuRzv
eKTTzlxAE2WlBl/ubDYcttsAIvE41ve1YaS45DmF3sjeKXEdi4wTjn2EkaUeIGKU73ao+DT9I1Dj
F+GANu/53gzG4Hj/SC4gjnT2A1wxVNGBLznPeO2QSYJji52UZcAqZ+bDW76i1Gr9j9Xu7LVgFf8N
LDRxu4cvfLnBsU7mxEXZxEKckKjPFn1jh57qtddl1gzmcds7vZmYWd85WsMn13ZDH+8EcavC3Qjg
GHZrAMf3zyDwLq07WjNIkKPvM/tnGnd384u9jUemkEYSCXhJjFv+6b0kKHbWxyXhdL1TRntwydpT
5koJCv97eTsb9BUlStfrTG5mK8ZYigZrI/aCeC35pXbevZMCxuSnXrMtcz2hzMBhga8Ywd9mMc8s
3E3Wn9yzGdNjpSw2LiSlKU+k9YneIAdypMr4shbjNCpDpDCv6JAQjwE3reTgptkTcwEq0wdAfxZB
8Z0QOaLZHCafcHG7C9dhb6gqu4IG9RVx4hcs6m08D/RZb6IRWaK2TTntIlq/EOhJo995qYOpSzr0
sBWMmxCXSqXyb/YgZK4QQE8gYvpHYusaRVUhrsfvRDJEejJlRlMY5DMatwI/FQ20wnHL22hQjHCd
J42Mr9MkrkaWuev/hHx9TvsKg1IZCpJ3Hsz1t/P1EfT5II7rjFzbjAZZmhWTWjuDLqtRSFYrNxSw
BWJFUDyFM6egjTYDP0xyU9RE96Clqto5CaLQOEW1ub7KxYyN7TpuncGS+BeOGyccud/CP9qHvi1E
xx9E2TJCQp1Kvrdcmi2l21yO4qx10Bo2qP9J9MNaoNlchJurnBzG2LUY432oYlUEEmsmFLS9wbAy
6BHC/FncZJMwELrXN6iX26WOSuYGyoRSGMvqUJZXVLc259uCQ5CXTSg0v8JXTlPaEwHbehdIVwbe
VfQtrnKmYNlmA27PAElm36Dd0PwjPApNvd3P6Cb/bQe/OLvT0+BAB2Gd+Ok2MafzYgzmesJj5ZHh
x9kPNjVwXzVzsgbd1HP59luVEfZCcLTZzSlB3rOgPjDunCiSLk2rlwx4HyDFvntGha9/qrHgRp5E
h/vDEzHNUp7pyWruJiMcMtHB6S2u878/JOb2pkR7m3jqorNSNmT+FdCvab/329mQOLRYbkoVqSfq
9Ds/1BYmJvonjlLeu/N3lLzz3zF4xGjwNnJa5qfKNC8EDewIuGW0Gf8BmygT0n6h8yOtZNp9qmjT
GldieIv74PzkJ6kYubJOPlZfYCXC5Akd1U2ZuUOAVIL8thSDtuFKiKpOfjNyPwOqTeMwbdo95TR3
Gs3hBmlyHUV5b8HwbfqxunXyqE9FkG5z+Nn4S06cXXcupLt/sLbeWH28vD7POtHidoJ2WTgamqtp
crVtD3ACBRgf/JxjrWe+k+8o0193KnoYP4w26lgD7gyM0yrfj/Trwv+unCZFC67dg/9uhQLNyCnQ
JrXBkKExYhU5nEGFVGQwjBzHvUi04wh4yczI6pSCxTwnf1R4xmUlENORO3Q+lNVIraB/rvcGZIep
OmrkSaTp2FoAWyl7z066SIiMTEF0w9dN9rVUL6Pqg22ytEzrPEy7alkp0fVv/tdHF49eKEXXWvgF
ioPHSANsNiCPghsgDC6ML13tyjtT26giawzZp6PJlGA80yUyLzUOTrGygPW3xgYwaGEiEWKByE5h
0+OhC3R04GUKg28tVJYVYGtlWj5hctEuMPdhg9OnomOa0S3aDHl5BXe+wlM0ZFhrPIFuva83eEu/
ZmGat7knbebshWHBRWwJXrMLCqXKal7WfQUW4OJN2UePk5mqnrfcVmR/zoq3BtCqE8DTTRgf8qZ4
uCh1NDLS3wIuPgwXvlK7hW1gfUzsI9T78j+Wh7rCJQUtKXtOrEdJlbVzsEgb9SJ1R2a4wgGKlnaw
yhqpG0+VdPEWgbPdws/QrRIjs9Qi5vLjeXN5jf0S3BgvML1BGPDpLDbS7l7yOKJ/kpmyyzgTCCgr
grPGLy6MbH0ZOJk2F3i2eRi6x6vlv0d1qnVZPCFRjEg5u2ijyJbUjGARk4mJWoZ5NhFLteBjRmAQ
0alufLHFLBIsxHkR9TSW1yfcqnGaX2aqRWVBGY+da2N7XPwmW5Qk+ocv2KT4rTeS1+QLvn2ENYyO
p4J8CT9tfBXE5RceFVfuREPl7jFDpuQc/y8XOlXKDi2sGzH/lBdQ3qj78twP4usMW5HUmQH8jbgJ
lr3gULZGUqLvUuR0yhEvHkNu1GRmALkBE5KJqqbQxKpDT2HqFTmoVMVybo9eFKlBBRwcSUzfUsRO
iW1paKWyeXysmW9puLNiqvYJuNyZ9RrYsY8k74ZSD/3p/zh582as/ctjMXlKHOHnoVgDF7nOh7An
zjxpOFNJUVBbz29SoEMhljMX5jxZYLFq0SZu/Znxlfo/TNxQqgTP154IfOdPifjYPjWlkvflOe8W
dR/t0FAcXhfgpLtzTkIICsp/hZ7Mpmh+6Jbfyd2tQ9PRJInMbShjWZ2pwaqh9yAMn6i/dMfU5RS4
Y5CIDY11tRbj96FvMG5tGWHxyxy1XPn21TxxwSgtzZvWzkDAibiI+d/FoBAD8jTKU4ZJspchfN08
UKYa7IvHcLBE9Lj2paKTndQIKgjpqM9jTdoIkLv9LHD4J+BYl5WCRpS1IDz1ps2aD3u4NLJrYezo
b57xM2EQcozZvKG/VzTvlTPRkjnIPL9ubbTRn8mQjWYKb8GpcsPFonsdyq5JhLgAT+fusI/QdrZG
d/fpLimcVgIsBxeQri3dRmfgvlg0x8ckMihpelFA0kclnc+iA7bPa9HrzhJKpTtBSjGvt4l63oUf
ywjzn64Y1B3wqUuLETsSup6+/qznra6bLCloHqayoXlZ6KY+qoizYaSGFx6jLT2WpUsdUk+7YQzp
BSObIXWMGwonkPYMdlLnC9NalSMxG2BiOFRaYJnvQAQiJ/T1IgL0BFy4toPEru4qweqB1bZxBW6E
aHooK0De8Yw+/y05UlzepXdbYAvo518FRXrD19rI7ngZZ62kJcygoltVqWtPCiHLDoh5TW0P3vxL
DxVEWVbQXizQQRyJ9lh9DA9L5f0ZnFQPVFSXXRd9A8c1DHzYv4oa2LrweyGPwglUB5gxVT2w95N1
umXaH4kptMSKbawkA7MODNPkpEGfEhmjqbSv8kuyQeRILAmOfX5KMRufMkqlqK2nlLbC9a18JRKi
5TvUall5QTLY0YsnDc0RyFEysgTPXBEW3OBMaDGAm1LLzNJ5cS1UgpcUFd77apCfvdsTQ3pwjCUd
DkDYl4Ju/82i9p0O8SpuVD9nBBxio/YU7vlAVFKbhZG2EPiH3Z0vZtJ5pBHwGXu7fFz7OW8slzUS
a4gLVwVYfHUkJeu2k7odV1I6J/XGoitYidIXIdEzR6MrLFLPR3Bkkj6bnuyUU2X2uxFLWn9/n1HB
axJZ+knBbq5uctYdx1C8dgC9pVemWxrSFvcW7SSMvFuWsY4WJC8tb2+f8yHy1siicalopBrsnwdA
W3G+4xG5DWkaahWLjTxKYc99s93X1AdqwU8VNVjkwoHaF+s9SgwfahAks7I4NemtBQrCFaYdpSof
rQGsK/QhTA6kqIBROwxWWR+ZeL+uqUhd4e9HBKdfkgwMEeqGBT2Xr84Ul+zyLOs+fDdoMoXuTkPG
wLOPWt4XcSRANuV+vCTzxFr2kT7y3TidI9oSNNdWQVVMJOBQvxxwXhjdxF4cLi8txvyBExzXcn+N
w6I5XOrttasMyG4pGiFoswxTUM9yAoEjobq3qg+FwbGez6c3kiNyh03AVeqYZMTk2ub7cUxkhy6P
H/p9kWqgQyUG50Dfg66w9yL6VA7vQxZ2nbAM6c2i5RN7K91AUOqtjZ/ZzR17JjB/89iFznTNQUvZ
or8qh3e3RZ0GFWpGlqJayX2pf1jOoin9Ti/S/PPBO/diX8tQBLE2H3l2abLgXL1hPisBUOyOY3ZN
KQHQgAWD2pGMuwCqjtItPHBNndCeXUc5wGNsKLj6EJFaQWUlsUn+P4hiSs8PlhZ0RMuG2kNAtWKp
3dQp1de2UHY5bHtlqRrgLcKR9B/4PT19d0fHCzpcWVXmtTFxWaIn6vS8Gs3b8J0js4gwEG3kVW++
KC5GlCipGitygd6ag9DtiNACUeTpeMtXk42s+4+HtxNYrHygHAMwfOUOXs6/dummOaysnL58lhjy
sl2wYgMFGYQkjGI0MUV0GIAY+dPsctxiQSBkkshNz4ItU7DSncUndWAW++K52vFn8sIJEZI6jhUQ
21rT4Qu2jyV5FnB90KiVgMHqtLisTsPTzuVnttLKSfTLrF7daQu4bDn4UgzlFCoupAJ/7v6yHwea
X7rir83ViNvXSnp9YWNOLUh5Uq95BAoXZ9WXENVGQoPwHcJvoLzBd8si/093tIcUMD+/yRP5Mx6L
Tpf12qEMLy8EYGvcd02oB+Bdfaoh2xaV8uCqmlB8Z4KfYcOkNTVorj5EQuzjvDeIVD6X7vfPIolX
WEYsfdv8GXQxkxVO6o4G1B272ez+G5eKYXerYb83jqn/A2VA4DZA5izxb8zkJEYX+PdvovN+ednc
guVwcmyXq6FnvNhXR7BTco8z4nklHW69fc+YxKxAKGUvSqaxKQBWW1v0/lTx4p8DqcUtocyBwTl1
ZnKfappzol/GJufro6A6y4xtRxkLDz+YOnJTa+OuUDWQ0dTiujzGR6LJjQXHHocEa5Q/Mjx0X/Q5
QGevFhgz/c6g05GE8GdzwAnHshrp/4ayKcXAZLbFKHuTIUx+gcItTaVP8kRV/CutXWuECgEDABbC
UEBAWcZynLiiwmV6zpudpGaf554m1yjq4kBw1PGR3J1gTneOYYG0URRwsR/9W7O99Q9yCwEiqdLN
BXF36sGmNB+vrm8lbirlHeSDRgrXbuvDWrhh/2FzNa6QqVIKWzh45XZY2heFPEU3phDSLMUleF+z
Uf5gisNmSXBzFVq6omuqav5FUexdCsJ0ZIRcFb0LFubnm5CqZFDt+uAjc1R1AyMblPsPgsyzKOxe
Rg9j28xBG/yGx0CQHLFWUjTVOa4aC+Y6QjGbVzyvNz3u27ABblKo1b9vaooQS0+4uGHO4EhZQULB
vI7ePexRY4Sl8ZojkbKBjVuMSjOPznKxSk7bgKpOIsJQKGSEU5iM+/RnRZNZLPJSWbqR9IGyPaDx
Oet6Khi/Gl6OOfX4jrRYQbOTNWuFKc2axYCa7ReXqaJqQoDorxGocQMGrnQ0C1/moPb42+7/pUh6
HDt9xVwQIRE2TaUTEir0m25nBryGJB6B0Lye/l+Torh0l1bZ1nJv2EJVf7jWbH+5KN5SDcg5uWkg
5fyT57tG6wB6U9+nv9Qmkg1mJlKIJgHaxxYoN1EErFGfskVggqFeKB6nLXCxPPNFM/WNCE9q/nYc
Pb6q8bwiXC8j8UAOH4Eh1hwK3FicmoVF8kKU6e8KePOEDzoWi6/MCY0VzTg3TG0e7mRCRlmaY/r6
hCz4Qk6kGFI5JdlhtM6QI9fTNZXLa0bdNltkyn3t+Sai2xzBYEHD1TshmWuBFrOBcY053m03C4L5
+zMT3QZQfPKABQAQPQytrhI4UOkj/lWd/xNqkACtNeYIFIZZ2qcWIHHbRQxdoek/6mO8Xog9S3Fz
YyO5nGP3TkeGXkgym0ps0S4W4Fwzn1YL/yX6X6rJSyIwFtke0W/eJFJ+ywYYMTML2bs+gG8KW2xj
3lvKq+d1VBzSAx6IkWWYLt88Ajvi1skoghqfI0XWK9gfnjd6a7eC6Aw64qx8ldwoxzkkwgIX4MtU
reb9bSGP8sj9QL828NCrSQbyHRBpTsOv2wbdRDgqdxo9BfAMfDziJwwRj3lFj9wxpQG5vcyp2qWF
Nia00lwUkeHswPliKYMNFjONHYYkjFycw0WNCR03pulZuoDYQPGBi+sl66XlkBVb+EcpZJW3cN4f
9fYNlT29oW0J84VtwClSMQCwH3fzBTLlkr5h6SYnCdp1+4SPLwx1ZEu0NGqax/lQNAd9z/3pPcaJ
O4K13BcFilrDMEP+lVvUtPNlX/QWjGHSPYhWBa2mv+QJ3MblzFDMzH689KOXc4vCybR2SvH2X9rG
V3efRAJRVpb5DF/xYT0lLl3IuI6AQnNl8UvxtBj4LIcoZcuYmvyO9Kbqtlw5MAgFbBLLG2IR6m3U
8g96dQWPUVlhPu5P5e+61rLiF0dwAC9hHYQ468jKI2hZWe7/VgHd8Gt+S3p6eTz5ONSL0BbWsBy6
ZPmUNyNcVenq/aJc53o155zJ7MYUbC4OVCtLpJv9+GQApGYgSRI4LJl+yO0aHu/L7HKN7XdDSv9+
vB1gl0Ygc9eltLRgOZUvy7YVukYahnYr93PfvG1aAxa1JunOCpqcUW7TxTn1W02SpH5FBF3hJPla
TGpI2qTdfAUwwU2bboTiYdtRpa+lJ86p+hN3KH6KRG5fq915/sBrqDG2nj7rjhr3W0F2TMpt0ZnU
SZ3TR488LLo9wOVwrUTbo2M+dzyDNAD2Kt2Ki3Zcy9Hwq6sOeSf3ksktolx78LPWoKydPbcWPAL7
XIenM+KZd5wLPSMAEPy3ELZdRqwwr67917DoXHm7l95Mm8AxEuqfKUC15IauGYNr4D7UYLzdHxr2
X3Kgg15epfSN8JpoUAPcaXkXUibVkb+UmRYUqMdTi/q2TZpKgLo6WA+DrLlzjq850x+/xzh8Mswp
/UI3VlmKu70c9T4C+AxuicvYzTtMJWdlaB9UzuEBJqOCYQau+Hit5HUzapSbKFq+2JE11YIRqQ+x
293T4AVKogPjZqbdga7+HbEFBDaOrJh3bIVFExgSFSYjsdXckadd3rz2HZJDYKoeU1KYIN1K7XMV
mDEwfLKf1xet3Nbxe2KoQXUTaxkbpOGnEGlR4irr8IJmlU8UAdXrKyo4ozIJIyarZVXZiHT88p48
SDsbN28F4AXw7Ru9BTMOa1u24kN3ebAUcnVn/UpIhGyA4CC+BBvwT2bc8Vi6RJeORnQ6AH+H4A9m
n6xJ/R2KEajMkZCBVzbizYcFJs5sZ92au0qLCObSMe9C9QJ7t7bdO9OXzN8S+nimbdKYkwjKKeWW
Yd3snEY6cys6+ajaszEaOrc7D/zydXi1kWh/qwHULkCBNpgjCcutLNKHp5n3VM4arCML5zk22igt
uNaYN7rq4uxZxQUqgl+JKRNZnNYDaTdbtocwY2jbEWM0tonhEQ8uJC6mb+GiAFkfRQNV5+7TQshG
cvkx0M9XgsllwycH3P5c4CidC6HfZxaeBPPuhPKIBje4J4aFC9fio1j0cN3MUpdwtgdcRxCqM63m
/UfFyTApDYkUSqHEryK/cCa5+morRm0zBlZI9b8YrjF5xKjQ4I5Mp0CG58wvKP2vfzO8/VEkf06w
T8DugkMjJsIFkYK0Cp9siyam8JrfwSnUPdwt2/4/f+iWNRhngi9vFDyqexU5UupbUjej7owo+RaZ
ffoD4VC/suw9oCUCM2abyFfR92gaOvZi7C5168sf1tiXPnMFxqhQkkhkrgHFzKVdUkvAmV6ejUxL
Y+UJkCGVHcwD9UgdTfQZQkQckvT9G9ID3lRO7X06jsWOz4gfTyPJT7E1OuXJipAuTSDx4KD7mRhC
t4reRlPe1NTsAP6v4nFSIq6tv1jMTJ/J5AICQI644Uk9URKjz3SHNPGr7B0ZmE43zjYS+fF2Kndu
LkzIET8MJfnnkpaVF4/9zKrhY3tPXFwLYBBYHm5bJJOzfVWqsLAJuw2TQd9Cds3hF2ATGWVmaeN2
XyeWWPa1uOqigIJXXqWgCj0xVqsySS/I/ETwxVhGn76XoT6wfU09zbAzkoz4VQV2BjUuh5pIeFwj
cvuGuOpmXQVX47ILJbtpbHk2kgOXxLRBLtDEAIKg74f82r04XPWhCOVZi6Wrg5fXo4ZA1CTbCQYW
spOlkpUsFi9TFsoctchKVZ2gnC3be3sJCmjAURWZaEVTJhAdeUZFFmCVn9ymjDAK3xWF1NlOQ9kC
d/aXqSFmPDpnrLGw1wlnFW3mPDPBD+UoVkUb6UyDkCLEs+p9GU4dV4EE4RpqYlBSf0oDp3s5RoXV
Q5jJ0hwBpsvlGtyzxsreVmgFVj6IDPhSrbH4AFwYJ7m/RO3E2gp74iKuxeg26rwJ8dqW+y8ZD/hq
u93KcwhUQOW2fu8/f9r3NwVfmXyuh1vH/lOaqGI5wd5P3Q+9A5BfQ4kAJnMiQLsymX/jIEoEE7kI
IvmwBH35zhaBKvkq7+m5cxTB6CTknI3T+PeG+z99Vw0nQVcvuQCWWpZ2VsNoG6fKYc/vviYS3F3u
wfOJ5PnaWBbCGyOIuyunSKES+lmGKCApuLwOlmrQUWB3MDWQ2TwU3bkljFFt0jLb1+fkssopQcWx
IKsf/S1G2KVSz2biNnT7SFPXHXMnQdew0EMyheAdO0nPSlw9Fi/DbKODWltopNQjFGN+IieQSqf2
Zb+iJQ0Lx0pT9C2X950ZqDqshplyDBx1uWZ3I2+2waR9+CmrNxRASC0afvEsUklNbp6iK+thzTY4
nLHyD+X2p+94HuJnfSRIcieoj/yo8+WlZ0DySl/pXlK/VfRS+Q0T2PH5QJVlTqwprUi77nE4ymKC
K4oqwdyjbnhbJ00oEhx9XTQ/aC11xK97dDqyO0dBRW+rXUusj1kdJ/DF9eoFOZuEBzKXeCWz/bRQ
zmhWG/WtO4sZk3D78aK2TaSt9Cr4uKCkLGbjiVZ9GglYGjBWpyhX9XkphsAipwl3Oaglcha5J1ZS
A0h1Dw04Ybcz/pnZt/wi9aL7Udb7oj4GFgSdrR9Y+ZMZfGuCunJPiE9235hG+53eoCaT+qMfEFmF
1vzQnccXot8cn2RZFq0FBkKmx4/11fREsSUyKaP28bwkuYTILiX3V7UPeTH1yCe3PEapkmEL9zI5
LvDJke5c1jZUg8xS+8hC6cP0+Thnq5giEK0pM7zfaoLR3IGXlPNo4IetwHxnzMdlFzkdOH18KvGv
S+IhFiuqtfAzm7oM3mrlyw0rGVLSarUvK8WdqgPmS8xha0tL7Oa7Hk8e8VuWPq/UWUrH+5QeVz6i
5JP/hdBGB+RmLRe3HH3Y8ixo1Zra+GR7NCTnJucSMbyluatrB7bBo0/VNiCBXQ3s5MJB1CQBANb+
9MwS0wKNUhVB4ipn8LSewIZy7jCOuCwINlIhY2qYLtjYOWO7Fht7q0DbACqvFXJ+Rk0XYNqE+HBU
3jUneGR/FJ9Lks+IXpHgstKn4NCPAsRzyChq/m/rKDgJ+5SaG0imVd+aMc5fUrumIH5DT84/VeFz
2SyYnhSjbQI6GR9IUmH59pDiiEl+Qu7ajAhjNFG/e4ApDNsmsXbXyh7GEf18hImm/1wJPVVpRWl8
0u4XsLhW82EFhurT11HDD1ghkABD/VyCpWH3TeW13h1Ctwp0nMrJdsaqWeUVH2rclN3j4PCs3l0D
uODixB9y7NSuTTiDPeKNErZFe/DRfFWUGSY1j97gyNFhAjEClg2ISIp23MJqth/aTMhWwhZR+S6h
IdG3+5D4guHXdmKOeH41Of+Tqm4GmdEVntdozZO6/9/X5828Sd/RnsPLfwGGVdCYlaz047ZSEHUV
h26xoSqGVDTuHFcIcTxTVgWKuowNvlEoViSXRQsRGUmi38bEcCSV55dgrLoYkYtyVInL2jFH0VOa
VS7/4rrXivJ/MI+l1mN8DoZ9CNRJD8od4JobEGlkamL/tt3YQuNFSR1Ao6kO+YhzuMn9jkPQmM0r
AfPf0AZNcI0TVa6KjFeXmWjYf2zDy9n7QtnH0cv+YCNkei8iSApL03Klqv2XYBcIRJe59A0uP5+h
G0X+9eQyushGjsbX1KEe3LGjlZyVjWWX/8PfiU7LA4vYfgAYyIE+iQqOk9T2C/+zbsuiAzitnxdM
kQO2Ck9WJrriGIAUqT3UJVRoYzHjgcztMTDvxalhRSMO8Fae6WfFeUegtOVOscoWNtTcNs3W1Q8X
Y9FbcB4xXMLUMVx8fOneUHNfB12qKaPJQaKvHsiohtS06eRNTjhHkDUv+pFSaP0T2MSwKEXVA3qJ
AXm+X/OuakbmX3JJU+DIa3G6XsgjA5HCcLsKPkYGNBNrocKOg1l2lxPxu+mXKdrU6g3YLm6TPHda
75hqRj/UVjkwSxYM6ri9+sGxtmsQKRfBg9uyILw1CMVqr0vWq9Fkl7mZP/ia9DulogypmoIZy1In
OMHU2nbKHtUFDHeetc9Ma1c9qY3DJEftpniBe0cFgoOu6T6a/h7FWIoEmAr7E3+b9vJQ6CVlWUPF
IHxn/1kMgKfoF+Eox3hUOkbhzQOZykrrtAQTRe6KaBnkOorB2EIbOPJlNWab0feJ8x7RLf3g7nBN
upmpMnAtRcjzbIcZLIvJnClkl9Jj96eexon4t3UJMzalAeOXMUlcfaR/tozVEZovWc/JsoMJQKBR
t9nMKRmt3CL/L8Ef187AS0NhdprjtKpBkcpUwfDqUaruVN7uK+3V6qZCvV5qO2PorjsSf4/F9XOS
QcuR8AoRvyV7rt6OJlGJ7Fbl3pn2qK3jPBsbKLN0ODJJGQbukj7lDhY6eABSeOilAR1EPtX0m6uv
vLh6FighRcpoBnKjREOXe9a46LK0R9bK8AXl4TpEYUPO+qAsfrulEShZi9yaQVNmts1OvFaKRYO4
TcX08XL9KkpsV4uD7p5TVuwl1LMYaBjmE0Z3tNkbLD2Be7GKvTwP8EtwD/6Ld+0wYUn0OY0Xk3qC
NN5cjxSdtT0tyo7igC3KwjlZiAwJTdtAgmBr8g9TLA4efCr40OFdsRIQYEi/dL/d16NNpdJ3cVlx
H1SDfUBWGeHP5RmzU/S9aExtQSpRiv1q97P3L/OVWvO5sq4BHceXDpXd4LtqNCL4zLpb7R4IKzdS
VF3ehlvjOZ2jyf3/jjW1gucmkR6sfi4G97B4ssYlwgjG3ieTsH1TiDLEfXk18az7SacpHnupoFm2
FPLDdQ4Iy5faw37oQ/Lsgoah1AGdyFZ/U3/tvEFmwQ98Yo6U8AXkJ6P6jK2we7uIvh7g7NUyRgOg
Vz1mq9fRRnsnFLOIg3eeeLWEfOj/Te4SVsI3YAGkqJ3L+I6VERLkx7Zwt36o6wnJxj/8aEscY3JI
jJts1gMy6JfM4+lVa/QJoCSf3KrR1jbCcZNkfjMwtYPKYGhO387idp9PInS32H40mXEACJVQlhgh
Y2CupWt0dcve/JOPpIsckIk+Zv1wKQoK9U2ew6nfRxunhDJRCVa9BtJIkZmaMWDibm7mB7Q7mS5Q
/l0K7Cm6NN9bxlyyqH7vt5NkLdSC1cjnARjOWgPoxI/3ijXZj0HqRjeFEs9wA3XxE3AJ0WpyeFNh
AWbdfNIp0vqk4ln9jqNFJZk1olRWvyARwKgsk0evkbJXUmGW3DpFbRAEWHaod5eZuR7FXlLIOx2g
f18Tww5AY62sCCJjNXe2PLJYjfwhzCZN0j+HmwDubleK+fNo/wZy5DfGkoB8TRUnZfK09Zav9Rq9
kEECG1jT3Ct7+T+VwGmKNRNOB73Ru+FZaW6ojGv4gmFYUcPN45iVxhsdGMcoU/nJcwyXHlbZMNBB
PaVh/7fgQ8X9/CLJwKReR3MnvOgNugPx5JUhen/KF7Mlno2LTIUmsWrtfEvSB8iLhxrmPMjyy27M
8O4/4qQADXs1vgh7MUWqSZFLirTKpVCcKHxJVvZ9GGP+/HtLOVFYJU2HH+9P+n9nK531u4z0zAU5
XHysI1Y4qo5BYcgeQ1p6iP8k0btqWOPo8+b/ucvRmDjuJHpF83fEUAEyWW9TWrzah1eBtev2d7X0
g3ehV2Q6te5WbzxWBBqpCcaVWKBmm9VQCvT/7emYmhR8FNogouhMkxYfH22tIxpm1R5AWbZ2BzRi
MnoT2ed5DZYdpnihz+6PDon6TBzxmlejjZVvIBYetH60W2NfsyWnmK1Cfrc32eYTbjXJoVqvzJg/
OrkrWzJ2ixao/t0O3guugt0kH3yPx/UAEZbgHL3frjjBVaKXyi1rAHnUzEMo8N/e1ZkHZgmgDvqY
JEj2bsjfr6lvAunWfor7MiB2xb23WVxyQ44lJkGibzpaOjRo4rHXiRoQNtwLGsMwWrqzQqXR63zn
wtl1yK9OTH06HBzl9V5mGjbTi0dt85TzAOgquyAqUAINCkETWFNBwqB8rJ0ZIlXLz++RtzxgvRqa
HLefJAH0NnPm6D/QXVRArnGK0j+TmcVf+30Ho8MOi0rRlbgu4qlBGMYZuepJ51me9eFmHRd/qWc2
m4CRG7KTFhLDu20Jp5Nfykl3Lso7ibXa1zk0+zGavV8LU1vZSsJ6H1E5OWF563cdj2gdgUv+IubT
yDU8FmLtG0ubDZfS8vOZkfLEhJmO5/1KevPTsKFvtKvEZY+tU+8yMaoOSV6hUmKZx/yS5wQU9JU2
AsbGgiUSvgs7upI8qo/fDfbYrhduOuF2k2bkMtt9PDmFleXvEeQG/ZBDgoYgok69UPBtA6SAUZXn
DpU4jHGB2ieag9Z8oamDhqPZYtfk6Sx+QgXL4CrBXYroLht9oBGhnkf26mv2Z+EaFrYFUZhyxwYH
vgI0uc+o5WFaIUXCo4do447btO35Nhun5m+10vNbxwxEOAkJi3Ljpo31D1kdXI0mN101rFmpITYm
g7pW4qSXCnpPv1nELSvyQv6zmQXA56RyDIFsVZNr6tYcR1Z6KMxlF61vO/lo1pmlEBvuJUA5ZZWu
U61NXX17/ZAvLnKCGymU52t6MwqeNWTz5g77Z4UFzY3PzSvW+a47deWF1v6jLuAcJKgQ21n8JrQW
iZzuxXkFSO0rMjtY9HfzLRgiqM9zmc9hBCon/NuAYkkDWDpiXt7D3txMGMtk4MmV+jFiN9jIQxb1
yASolTY8v/ijQ4atg7yl7+vgs8UKikQCe0808hTcqNnzS4Ch9UVxM6BBbAhCdws9FY5uCdLJ6Uwz
rmWTXBaxtDFLVrQYVzlA63Jy6tzHQyaNfLbMepcyMXw/WO9qva38MLuBGanIs8h1LaKuhqP42Om/
VzUh0/y60+ui50Z6H0JBJBlIem6b1uZLZLY472vlq080vHQt4rTw7XCjzJV0/B9d3TX/eesyw54n
d1V48MSo3a5KTHc41NRDLAyiRA1Nafc1jvgfxvczpvEXOcVvS7mB5Ff+81eWM02OlEUsZE/nOgJN
PugbZ8JEpISYwsgodWQne3eN7bay74i7J5xiTBamWt1etTBdI3rXM1vChXQwifN+pWahjl9Bkk+h
YB9Ka1n9qaKLUku42dgGleR0wbDJNsJrn6OmQW8tNErwzdKzXRADYQBdRqJ4HR0tzRm6bqhoST2y
mT4JR6JhsAQOirD8aAaU7+yDGLCr6mYms5n6uOu4y6z7bP/JIQs5/AgS3gP2h2vTtqNxj38dVr6b
THcEe+zO8+Ps/n1Eo69OCl//8ZckA2xLsMJ1cU0iPCa4epRTqvbFpx7oVbVG6QrkTlA+jaI3I5zJ
XDx6lGQOyhHzdJrZcpMbINgVE5sRHCb8IKFuduUiRHTYJscDFGYkFeTP+4kqgFJm+FXynY3ryXC6
un52qzRkCvtt4TKAr1ZAbyUUqDgu7v/r9xvgsYuAKBSC9iV7/+qRMNWXgWI422llaXykdfAq2ZdG
2zaYhdLPdbkldD0u2V6ZzQHokBUdH/BqGc/yiQ6IxNVnXsLsLQ1J4S2oigmDOFY4s1/Lb+eQq6PV
eQE0p23SzFxeaioUi4AJ3djvinxYG2ER0M6wmDQgyfcoPykETnjS3wsxDirS03t7JjR0qvYAFgMY
Q+zmCI1nDbqXAyQuBIaZcu7TgsN7mRh2QhHMh06YD/lk//LXIU+1yfwIBzr0/JDvtnOSoJ6LrC6j
9bq2/kOzK/+K2qB4yJf9Sl1gGzNSTqwO7FMIsrmCeGGwzvRtvXPIXER+2RiorgdbQc9ayQTwFDU3
l5TcqX9cOX73wihNTDtPqCGZXBVjhtcawzboalWADQj/qf6nl/LdFfW+27PDiAKoswhoMS5vOtHJ
KP4bAuow8pcrSNCbRyyabYD0r+foVOq3J+lnDk0FQ264gRwUAlkk25MUAueHqOK12JbiorAjPq9G
NQhLQbPgE74aLDLGdbtioYtdr/7tlS1PLPOMNvuhzTupwuId+EmYznY9JGgustA9N4siuYSnxII3
Em8kEx8byB7Z+sQEqLq2zjPZx4g1guA7HRSD8C+zu47B2OnstHQLwSUqSxZDfWEYC719qI2Kmg6I
tdXOUltee8h9mGJRERWRCaGPwHwKbyGXLB9URyjc2vNsXFDxaEaNUsoFFpWSGvC4+Ui0x+8JDe22
cw+xvH0244zWPneLn0cDzcVDNEp1C93pFNzZ9jsyqvg3J19+ZRtG+hmGbUJgYHw0tEkY6IyBRBoK
W5hLfGquvet3jn2qAjI5/O8+6g8cH+QHg4lZ7JtqxoTjx2+VpxAkUVX+kuhN+B/MP4T0A8/UfBAH
pLyBJnCo3g6UogiHJXOvj9uyVO9AowUljNaYa7poYzJS9yWBzY3rH2QlDPuvQ46fsp818tXwMU7E
2By6cm5SGixL1zsNUdInEEydvAUSXIPQ2aOCs6jZ7rzyWA5Qg9AErGOBjIvYIyl5Tgq1gkjpA+Y0
DiyQ3hSMA6Q2OIK6pMwmMdOMdHzUy5W7mAWQXAhX8FN1umXJc6r/4pZO3BzlvjWQrBx0Br7D5Hyp
3pRF+FKA+fu4mFKWi6Wv4BGtzuYXn9DDXJQ8EbQEiqGEiVh3+SRb2u+0wsCnd1iRd1zxodlkLVR6
5pBFqLjr0iyG9qb8Oy++JbTA8Iig7Vk0X36Cue8nErYDwa2JTCIsprpYLawUHzYumkUpZeLg9g1V
PZ1Y1lBZHV5Yrc6DZ3poaN7i/cJLm67gSWX8hQH4hjPkak2Vsip0GtzY74GR/NiIpuWZwoHoyHFY
9ZZ+bpQ8yq6hvju/ox8SaYzmfUoWfiqVCy6SCD0VMS9hS8JpOxqI5pqVfI61lFQc7DbGHPrXwttN
o6TkEaFe2fKpwrDylt9+rVC6x/HsEC2TQtkO35cmub6KuE1FonOQD7BErVeLo/l0TBJEm+/E9zCp
RCMUSavspxIlLi0fvrkeErdmucxVc7228X5gSVUvvMjXQOyLxEwU8aELkVCXVaT9TSixSWB6oBfo
LSPftCxaDiWlDtumadE508E4yfrvXWmzVsLJF5KrLCA/Js5cDBxnc8JQwhFlqn2SFVXSEZXt+4nd
5ApQkwzkrEyfSNB53cNNaUwLxfvH064o8lLojSvhElNA2OdZNAZNd0tmVbaXn/q49gZJOullE8L1
+8q4pZJPcpHdVnvcCtg84AHgISpEdK2UshJuUY2zy8n+Qdhm4Q3W/j8fFT0i7zKcKWn4Pzg6dEaB
hPzLTghot4JOII4jmCvDmwUrQwJUgQpgw3ViyLlgnWnS89jXBIUUQY4V0+IHtpZf8l/1xDo+CTKY
JfDVhq2TUxDu1QPRmDDff/aCUCl4/YUfxi3uhPhDsJtjKIbouFMhvargh3Z96uaB+sN4Sq07Ci+y
qTDrzmlaeaR8UrIs/OAfITWSUK1M7No2lHjzk8r13A1JI4JZ6VtwQxF6mCqIEbxQ43IHTbmz46L0
0nkSwAtHz2GbfisvMCSh1iJyS3WM9oyF0R11jxA3ENL1FGkzB3VwSyzBhy/Z0SR5B+J4HBuNlqt/
AIAipZPYAl+aNOUCxxU1hr92CpmZrV1ebay1cEngTtG4BvGJ1EHyjdBpE3EcsGa2hF/JlQE4nPAs
M/E6UQI/1729aCdlr1hESrZ3s5ojHgKP7KlYpt5YkhvYfFHi/Az+CZQUTvfqgAm6fx/zn3+P6XT4
gtVvwoUecXDcdPAsk1eqehRXwwaD/7/UbhncYtVnSkIOGy7GJW7Dockbeo9J9+Pb/biDfS/T+f4d
RnjdMu6iInyry0o8dH5PYMqItViy9Yb1GRPIC1Vb7p/BYsypHN7WUbs9h8BTouxtkGs4kQyAQjKp
qwyy21ZZTF8VZpxcdmHluas3PtviWXdYL7sLFCDtQJNoBlDpu5M7UibqGAlSNo5x1xuEgqjN1Cr+
tB+ZvydajFGuMngXjU5P6QaXebAn5UEq7xchqhAKH3XxKPZcT4kUspnzMlgVCmWxz4r2GF4DoVXT
T60E1TyrIN1GLrnox45wUbCfMxyEryKCaaIpNZRQ3MV6Zfdb38avAIiwCaJP3w/xAm5LGqPviqlq
phXxkydjyiFoKcrBS+e8UmckJZm7ruULP2Nhb+ZpQhStdUjV3Jz1PTGQQKQe4HSSz5dpyCZucRhk
VZuXelgJj5o2r3N7SME8vQtunstW/c6vj7kcNx6sLtKZcDGkg0iybUh3hRKzenvR6eWc+6OmcQfw
Rc5mNxV8DG3gvDy6a4wYC5rF+umm/hlucOu8iaThBok07JpvZ3nSG9xuaH9VNjxoPW/P6FDTcGQV
KLURpNAqtdcKv16vL72QL3I7RXHVnfkYb98z0cFh3b0Cv5fHNTHyVkWrt0jffuObRa+R9P5cyZUt
cjbGVaNJXN9ZMN4fZaeDdiEDPhTpL6khMp1med0KKsi/Hay4EFUw56wWmiy7PY6zO5c2zzcNbsQr
TcdyfBqV27pHRb2U69jZqhPbWnuQbt11bt6zaMzpEzle0CiK2PjOMIXfdl5mlM252POuCoCCy+l7
rR8a7MGvWS/xKn2h33qGATaffLd35nqAYXDc+oV88ubFysV4LiPiz0pMzlCmvTtSimLpCNgDiDJC
vroaNGKvBCFdrm9CAdvA4YhMt5FEZ5Xoj9m3GcBRB2WEifPEq6XyWM80IC7WPpu+r0+UDPIagH3y
wzLDInT9P1REPjp4lzUcmOQuw21tQHMxRxr+LG0YWfx1xkac+d9D4xemZvJ087k4De471a+Uj3mJ
YDlthZSEqozAs9Tkno05f4ciOvuIgvqFfTZGSWrtatwHp+jdGnIm2je6pquB9wCWOtrN+JGPpsTh
WjkGXTYtrUPYVom0WbqZ0n/EKTvuUG6rTlmb40yuk/yJaA814fKw5V6EWrBeEcRSgnJOTL47beI7
UCHyOOQkmqWAjon5U4K92JowssZJ9qHCdMmlSRDHD2vlF+dj9eUoBMdCll82D2yodWXlOLh5BcYx
NazT0l+h0ng02oDWSY1zSQDRHE6lYlsbvxEyCVRuGYMxFl8zF6YmezKJqZCIYI3coNmbUqIt+djl
PbcaPnbnBT4meBzGGliLBPy55r4fhMvk6qqTuVlCkbRz4utdSmLoj15nL3lZWqnCQxjLBxHEgEp8
t5tc87JcICuDrvW7GkoAhuQo+hfWKnZn6Rt9I6F+12xiY4SDEy39gQFIKij/KO9nrnVo6EWvviZ1
IDkxN7gUx7KrhmYrXhsEQ5igVlmY19rXcZdZgETl33yBgfO4SyEtTw48QjEfjslqMiTplEromyp6
bktmIaQoca50Rfj8mOjgy/Kr/nAGpwH5miv65nPC9237xz6zSHIo1cNRZ4Q4IvlASJtm6jeH2dEM
gOG6oYEY7g0XRR1iyoqpmK414/q3EuwoKeUdTI3T0DQLkKFcSj02wDvWAYgLH2wPC0q+rz/ZTlAo
HuvdG5ctiNZOH0HL3iqHhuBsDLH8CWu/pMoHdbcKH54X5UgKw+i0ubBw1rFVj8nGjJMxpkrBHnV7
AU5wyfN1lO8o+zRn0ZglccdAgtv5ans++G9/eo3AKNCNum51lmz5ROG0zsqw+kuWSy7VHW7Z+Mia
v/Wiw93F9yYPHT2jeg//XpbkvHmw6YDar4F8WGihJB8QBVdxL8rjPJofL2kpx46/5b23PZSYff4j
K0rLKUj4dqQ/7yiY3LPfAbmgLxvXsehJaufPKOvR6rOR8DuP8pR47jLbHmVD+dSzqVDo+jNOYkJj
/vJ/SmmssJFwzpqEGg+NSGNCZTCvA2q166VlExronyJybmSu7i3OpwfVP8EZryn5TvgLgXc/XOsg
UOuEhJUZGobKlltmqmv2iQfvKRpCZznomevvjwnHj/sCmTod1r6pEm/Kw5smePTlAhBtNJ0joF0C
1QTp5qnR1ZrdeI81cR01BCz4Jj2cikdWgUnNWofC1sKzPyyuC1PMn2uyWd7jtgkD4NXaa9N2h1Bd
H1erfwWkx20Pu3/E3wZQmHJ2gcYk46qAqRkW0WChmDdxdNoO70XkS6T3za9JGKYmfKMg0zeWgSje
iJmt7L8JXbtOQmD6C8IXcr1OyMAte/Ql3+ak4yl069V8r+6gwnL23j8hqC2Qo07AkOmLhXAxExTt
vQrmUBpwE2/E2eTAavQ3Zi5nQWxYa375QEm5spaYsEmluoGiwWgJz37iTlfApuRQ344jp4Ic9EP8
i0CPhRcm+vDjd1TJ0vRaItGjkBzf+j2+N1NOj8MJSnR1hsRDhmIyC7WK4P6YFI91r3V1sQa/IDeq
eI2QkfbEQv4cY0ZWAQNfil/k2FU6otKZPu5UyHjmvc7I1wvVyYm2Y8xqJVTM6USFOLErIODglyIq
C5Ey0wh7B9CfjHCTKs1Ef7b+dKyzkkbNW9m+L7odwZNbcn+TL4g516Q8klQZhfqWw2zMCm9ON9RX
zcXemzP9ZooY0fF/q5ykBhdY0SyAa8g7siGdacASJipcjwxPl4iKbNbgsGkapQIB5SpxNGNN14La
iQuzbgEZaQ132JMWVM+eRptM2U9tsGrA9C0aA7WfC5zieQt3CACSA4HVJuw+78NNHyMGL9qeJRlO
MlTr731KymzyRVstIuikt93hHYzZNFYr3/W0UkEKyHZr1owLRUgmAD1T4BHMk1tWe8Mv1fbt6iYD
snJS0pSMvoW7OvAU7ssk9vMbXgX4Qjb3WauksObB7CQV43P2omgjAmoPNIfOVv9uZRPgTLuBronO
3jR0jCfeRjuFEyWfoUGlM0DrvXPXxCKYgayaxdNB0RPXj8BRsjD9qmg33vC9jBxDRUgDfC9Z+jwZ
6Q5jluRUSPcdakJGBwhvzJ1A4SvwfBgn6UPkrWYG2vB9fRWf1z5HQSKPYghIRCllV1JDwcU45GQ4
79KxatAKx6LmoqeFwnxzyFBUJR7GSCm8FDLUdPZQ1qIMBo3wIQcEtHlhl+HAj59EeR40/1d5IDzJ
dcNYcDCzXncpNGv8om1i9VRtjM0BItUcLCtZKkDZe9S7DpMCPWUiCJwERR6y718GmiuUkCSie9hk
Ip6gCDdkh3olKt+D+oADduP4SLjeDPy47lBVE5LBobX59di3FfE6yDeyxTDcotPp72RQwm+Xs8Au
vpuYiYfZB1W9g65TTvXto9m7/6/K8nFQZsBbDPtc97bosk+zgCY7F+UrhGX6VYXs8JTwcAWR6ARu
TyX0Hy1NZk6JAWXwlmyIhvzy8Vm0onrrPYRrx690CObgjnkbRJ0wezauebOFJb3I8pP5l/cJmQWT
X6LcIRnlmLar5xhKO9Yuo9hDZKmAWydWgm1qsWSNq0fI3PkRz7tpbYCgoXzWxhy2UKB8cTj19j7T
l8a2r8ULV8rID1ljgs8WGkqtTObJx99ZVlh1cbQAUdb02wEBAwr8JCE8688dz+cqgamvfVgZgi26
PeFPywQv20pzqOAO5GQW/zgQNv1MgVmFCYSno+0qbbfFpN3koP2Jz9da8ykiW4Z/jzMh4oTDz8Ww
YBoU1woVNCBEgA6ZYAYP5OxYtPqoNB34AcuyKxQWAOYcGN/G5ZiLdM9bLamVnD1l6rzDzGurDu0W
Vr28ymUeJIE/wdPqTKgaJkkfPDmM85itrd7DUgKF95jri4n2ti1ugWQIBN/Ey1sVteFiXay6b1pT
OL6nbKwXDjXrkOzrGsVpDGnij0Fjlq+dnjJ9aJoDYQXN0fb24qKduT+DeVLtq21zIvsb3BxclHwo
zNYpJlDieAxcYsxXe2Y5YS0Sn/jK6CJRMyihv6Ca+uwau77P/a2LxbvQEfYKv1xbAe/Tl+YzZzNv
n/00LS4YuiVzjOG700MyU6TheIliSegvbwst56HIxlDtsnpg6bXk9IYBZnBqGDdQKzdxopDfE9qi
ILnm7sz632TbAn7/RkQBb2e4naXZsJ3WB+LRqk6+b3zLOTkl9zdR8+GSzKbbB+EMfSICmOOZ/+kq
edO5YKfHudUT6lHUDIpfQ+RRrMfaQ9MDWWMLOTobkXiZivFuy6xNPScpF1DgAdYu9BxtF6wSxuWp
hW1Mh9RnNtr8fBOy8kSYjwy1AqA5eXF5lLTzgMuT2qV9J8gx588g2+NjYxaBjcSAnHx+r0QdyFfU
MKb1tw7qIrSo6QULulN859E7Aouf/yz0Dn0BDkb1a0luZTZf2w8P7HK9JNpqJOw5EynfEyltRXb/
BYERLoetTuOUZGTcp2zDVEZHlm7UklEPyH0IFcz7MzlqdZRcQnlpuFA1+5b8DeJUMFQxnrotFM+f
y0eoQrb4i8SehKoBMPnt4AClglcjmSiZt3/47UM5lahdY1YAgzjCumsu3QhQlNyKS7aZfbauKhWt
mZrCUeIuHxOoaN/coGd5L438dMfw7WjCDoEaEgmDyhhL76hYW5+qB5NW5g3balAnBq/KV8N9K5bi
GQv9EKwZvpJ32HSwVeMr3daI7VsbzUWZHWPlGmY1m9OvI+1nSd+ZqzPsqcNr8tTLtzSTewuhr1Uo
g/OJlLBVeCi/Gl0hv4d64Lh2h+EaIpFz9sj7WE1M7zTir8QXcm6kAqPtT9nTKfI9A8VreKzRgZqW
8GOtjmH4AFH3maseiQj0PqOhmZIeRWXDhDJ1iDa1B1J6HAF42RMdkOQUeNFmWYmmkx8BTDoIeEhu
QDziGRWmgGMr4sk2qNNx4ULJjoEkZlz7FEAKOOmLTOG/KW0ClrOq4p5pbF3u7ND6Hg3tCiT6REB2
dwe68SkDl+/bd8D+JiihLVwLIKvELXrNEi6NTUPFvKnhtIspZPjqdrydToq18efzuJlHWgrMZzmV
7OMOw6mAmWiTxcW2DY9VM9fI8NCXDoJ8X0H5ibXGMJMMCCurXJOfWs5I+sTYRt8BU1Wh7hyKnvwH
skgQRV3Ta56/IqENlOhHUmyOJO9TCd/nZuXzw6T7wTCZzFRujNGi2xXmyQQUcrrPGIKJZegX8xHv
LXrQQcXDLbjqV5w3efUq/8WljcXKrLzYdOhz5mBZkfkT0K0VKfxmjSSkfc9zfU1yCBa8t3ovxuFM
50zvdw4I40gwNr26Y32i8kBW8nIPPxc+dbvAZ2IHuqTqN3eDKPupAf+KZVaSZsPAOlw2VUpxpfPo
rDX7tiMOwBMJJsJeT4/L/TWPA2X44jLLipvKYOaGv9XRFTQBTvARtObHz1BLSbMT9cLk/sBWoK+T
JyehZ5LD4XVzipck/JwO9i2eg5LXI65WHrvSsqUx8IPj73ZDLh9G5JeZxWwwMRhNmKkLJsPW86jP
aRQK4eNZrpUSliriBZzM/wj3W9D5bpvcOgDBX/XvNa0MfunUPCzxl5Iu9yIKQypWSdX6ZgPENLIO
jzb6SnDjTunjU054/crNPiqG3h6DrhLzZ2yIFGNhwS47qOhUky7sZoWJFGcivt1ts94GW+LaNiAU
t4gNZgxndFTgG9pPK41aL1/Ka8KvDBho5sTqfzYIhkA+/wBpppXPy6L0l49TdeP1tgCEdoFiRWo0
rRIEJAbt7CjvUgCGAfRyrRzod4rhX3MqDg+CzFLtZaM5ctJsMHz2d4/zMgw293zmIbvnR5BY3o5O
4E3RKgK/YQZLPS0KCdNqTqVBWhnwBAPmnJX14h0x7Lt4TG8YOBvRiMtJkVpKb3IoZnCoieCVg0ad
77T4ASmwzJ6H/nmmmQ6ra2eLL9Cw3KlF0HjpTadtW/NQMo1SzvFNK3CulUbEFcV/s9WbnrA+0V/q
6PCThvL3WL/lB4Lq8MidKrhWyNe7cHHdJHh82NL/4yq1Pdb7B/ImNq7hMX1CgNabXMeca2lPDfrd
EvOrZVPMT3pgIle1G+zDoSxKDKY2gMpP8sgVXcDsS1tR3VkZMco+popa0fOmQY8Lw4WRJXnIBguc
KhL/sFwUhgku8nIi+gypLxlh2o+o/IBFKgACeIS6sRSg0m7/A7AuxrrJ1UOCeKUjp40/eMN+hNpT
0QCJCT8EecoGxYVHVcj5B5cq6EskwJH2C3b3wlXYjOvelqbTxTaLpxCSLMEAhvpi3lE4S/rPNpBY
pHcR+klOSsbt38YOgAlXRGO/dcY5bLRnfkrkoZW03JKKDaeA8Zt2YW/0VzQQoPdJhoCuG6iApGUt
XxSNTepUQV+KV4eyRzkAxA0p5MKu+xn00PGrXLE8/1NR/iEq21PnFYGgL6cTWPb1aSMIMQ5oB8SH
LZzD083uw6cmbPsdvvMS1Plg2xjIz4Nw4M1ESSkm2BpmxBiXpDOHuBSTNJT+TVVpYJPiaEe1M+s4
6Ea2Guieapk2HNUGEld743Lwz4X9FDCsGDOj5pyQWX89GkSdUt5RLiQZZ/0JD3JjWfiUnvuzgRTf
ZrKauipbCa8C8I5bFFMZn5tUcZKGSxVHH28ZEnWQ9qKvv7RMg7OMNLliBVAwPVMnBt8yIWjfuLLd
4qKpKej7VuLh+Fd0hA9M74kq7aJ4x+f80E5KvMcoTwuo5kSb9MxuDSvKDuz8WnYxos+FcTXrzj/o
coOii6UApjCiuA6FKsV0gI4XvFXKr0RsWZ1LZmdWg6JKa2Zy12iHUaFrMaQ+D2LlpkP/OnaalnFN
WUuCbYQpeHlOPek3lXcdAWoTPIaUcoga465OaYkbGR9DhAjfhh5JSpnt3yaAP2UwWZQ5nglM4lWK
kq7x6YdloeJanIKJbs+ucp1cw4IU43G1RMAqFzu7FKyD4TT/x4Vu6oyuE2HsFLZGRuhvvW9mA+6T
YLE25Ic+XBFVDtooowK5V+2TNBQtOxsmdeYn6mgLRnMkg6f8b0VYv+fTTPwO7PbKS1f7UGJYki61
F5UExzVSXly/kR2c3g0KVn7W6vJup8oVA78rrSRXn8DZxLqC+vQrSvowUg/kW9Q23Zn1FtdHXqqQ
p/WWvIDsHt6BYPe7H/p+b/boBdinHRiO3kG6U3PlTzltVQxsQdSuOFRdvZvUVTZqtXCUKF4gSVZc
O/Jk5yC7GqpXLl7RzYZOGds+Dj7NoJuD2HdT4Fw5V+pSItU7slE88wfPLoIRbWUYG2pp64S39Q2x
GB6r3LQ6G1Q4fkugP5KwaxKQLCByVAa3zs0whdxYf34MdcCYneICkRNedpTMMW9CL/ficyElgRpy
djJlQwLPgMJ130vbcQt/JrWJFs1scjtDiqLV+s1mZnQ50io3WtYQUQdro/6uYjk3Dy7Fv7o6wGlH
4aaHpg6d3Dv3AxCMgm0dIrB6zOrrTXRaYRpJn5GhxPDg0Dv95rO5NEO/BbunMPMeJypdf/4zAyGE
GVGT+hMCeSBWsnmtrMbLrVRmRJId7vR/53RS3kM+lJBS0k9JBil/lIJTrXWT13+nSespj+nCpgYn
pFSEh/wgf0Jb0qu+bI5f7wONSQ6YbtBnNMpOGkfqtUHQk0wMZ0P+QUwTuAkSeXjHTZMJ73lSFcDn
HQ5gOPXN3r2K4sz6PCq0FR7ywZgkwjLVNkNP0JFmrm2fEdSQCcrw32STnuGbjXdm78dvrGTgERwA
K+OZf64WGeJUJEQdBJR5VJJEalBid3Eqm78EaTb7qKYUypHHrdoSKi4rTXzE8w1WbG6e3Uq9yS6S
p/Qv9lzrAf3+oJji+lRp6AGCC2OPnoo22GSfnLYtRFKN3A3cVD6OPaFfo+iC5vuk+wJ5LwZHjBN0
eWU+JU8EcpihcnErsbwc6Z8hyXIeh/s9qxYFtPgG4M7V1Ke6hVz8cNOs2WIdrp21AglnHEjZXo2Y
b0IAKgzIMqDgRWjSJm6L5SuqfjXI6wy2l6FSdPIRN69ElZH6PDarQ/rmGVnCzJ/NmdrHL7tfyXWy
Jv4V9ZKMxTe/Da36JVVHIwSqVqt9j2dLzGetHvcG4tfNkzasqkH31ibwae2WUEc2r39cIeqhBhKj
HVuOnt9yjRng0nxk5G9gXFAVA6h+cIsyQJiOoJ9H+rgQjo2BMwgaD76MiAbGsU1I26xv0U9yOoHy
b6DqkBpRAH3JrwHcMvvzlP56prkpoWV8eh1Cr7uu8pLoP4fCTRIQevHl55oz1V2Mkeh1aFxRAF4s
U/xxCeOExAh0v3KCAIesQ72wu2QIwWKM7HoHliQ47CWS6SrN5ETwfuU/52pW90dhYtsLXb+pXUrM
hTXohXQSIdZ9OuYyHTUh2UH3lGU9MxrwWf1zki5ZQeQASAolnSoLO/Vqf4ATG2DQB2pLCoHPOIie
qY3tByIok//tv03GxvuE4h9/IjofDJMfN4Yew2Pz0Hho5UVxK0NFB2OiB1Wmb6Khccs49EWfcu1d
Vi/5hs8J19FkJirVVYBqApjAqV3BCUDNBk45ijthb72FWxWzzlzDmS1m8InVrx2d93yHm/HQyU06
PvtWj6BCgvazI50Djrl9Y8KlMvH7WLE2C4wsXEGSY1mVm7Q/UlbelPq3KjihmpwaFVAQJbjvqWKP
tkzv6+98cmWF5DLiWbrrFcst0j2at5+ic4XP5sqgRr29/5/oVbrDObQ+YsYle4vHKkpj4RvMPFsf
bBvdOmIuqSuMqohVLHMYujT76IGHtheZ5bhbRz6U/+4ZSdmIGNw97n3aNqzZH8zOykPXY9OdUsH6
tR7n7s0VUPaJBmntbHX7agyT/Gm7BtKWXwzFbAEcdVw38n6EYo9iH83k1+y6hNB7yNSWI0O+pR7q
pU/aDKK37l0CK2FRrfKgLwUEnH3q0uVG+kq9oMh+Xpj3d6FJYlOqB6Lorl55Fs2S0K7vQWhMQ3dS
wTXD8a+8s7y061VTrZbeIDGUp7DHhB3GsQ3PehreuTooXzFEKSH0yJloZ14RJQXAiLcCcjICt5TZ
VkcmXpHvPcDXT8NStrMmDCFCHC3zbOy0PICaOLOiX5Eniq9Usio0dsfupJZnup1F+NLN93oN7dra
EOmrRYFlC6dG+ECXRlDeeKFWMpxbmCoaCvJccq5RVb3eVdLmZ4if0IqOsSwr1ba5/rYVcq1jY7OP
de9IbPLjSKCEJbRHYOGDIUndTNSNNftTK7Huo43t92sBWVu8oKS2Z8TVcaOSL5FyjGc44UHtuJmO
tkuN6gCxzq85SVixsybiuVmnnWmIRscFuW/MN0Zdt5IaGIlxKdlZ/5gj5YtrqzBXmYleQ2NxB/Sh
H2AqCsqfjhwTcMa30MSu7u2OV+R8zZ1yq8pBDRFzpLOdW0hdR/dxC0ZGkR+ZFwFLQeX58IiPJ9q4
CGnWTfhaz+f2O2rrefbvMsB79kvkZGUMyYeGGbndxxz5hV+3M/lqSDQgFC2qMHFwQuRIFKo9n6Tw
9DJvBhm4azUtorHb2CiXmKrrHPtx+wPEhSQkDQdwT2mwtzbfln5eSa/ZQ/RT9kYtZWDoyvB9Wmod
HcJn34hw98GsdyHd0zu3LlQT0u63SoeX5tSuK8XfBRCgibd1eYBCC3DP5WG5xdDKrofrlskq1r/w
oBTZqvqVBwtv/MOSVsd+8u4lobEkWRyTebTn27TIYaOD4CVYA6SZ2Y4YaunyNQBDFk2ormquz4+9
nwF+pb9ZL4imf9kHF/d4RbH/w3y0KQSdAoSHaWuB2vYu7gY5fxmKfwPMKJYhvNPNv0fWypCpSsR4
ZZ7DzP1GWWDfrSKM1NxntvmrCyJ994lfAIcXgLB1q9CcxemPmRlV1xBLlzYiNgZJC7qygAmFIQw/
dvIP6UAkTVo5/9HtkuTJ3rNVhDr09uGVK0Epes83gWi6ogw6Mo6gFV1jgR+J8y8WFnSEST9uArKQ
ix7xLtbs6G49OCEsuQt35qsyUh0MuL4dnZzsG8A3NKas262JmkzRdP1A2s/dRxPG6zCpx2lX118h
aYwxBDhYKu9wQfC77fP/uuOxcOVPvTD4TPks6VgRmuwIO/qkNyB+5PyQmg4einA8kTTN6mn5l7gx
wSTWW9e9UGRB9qB/Pk16W9yRapIWIDxyTmBgJCresxRDF4GD+4kT5onmddv90Ib0wzSbR6W22G0p
ykQdp5g8ok7SvogH2o2Cn9ohsN8esdKGbMXcMKXYNXUWAXUJCNlZ+uMqwKmecS85jnkMJKCV2+cU
+Ce8zuHOoI/NsIH/8K3ukrMWQkPBtLJQrVKrPNaKos4vr33KEPDN578Pk7UFhYkpbqwAV+kie5pz
ESaIBQN1QgHduXccsPZRkqRoDX26U+Ty2TOCItMMdk8vHXkN0XWGIRJmH338R+q/HQkaWVQufKSK
O00x8s6QgMMb0WVx5O3qwsg56zDC2qpkO2R0sMhgkHJn5l2H9EiPMcc//XOvblfPV2/ocuRssM0C
ve63u+2SlbktoEETEfHiQ2e/e/TAK3ycq1Tyl9dsqM93S2iVJm4SnXYm8dc8stXwrttMSHfc8dQ3
FtJbmdXvcKTA9k5v3nL12wSzuccHBcXPd+Z7UamhOgEiHAcNeA23aT86MRCgGwnOPB/GrX1QWWGx
lV9GjtsCvG+8C0RQRMHSbDRgPsNAb5UTaYEME8bEEMKEH4MlwNNf4Vs4y7Tjv5pVW1mqtOmcu1zo
YHMyYAKYQKvf75V/ax6pkbI9EUWzpvCA72p5r6Qs3zr7ffHIftq3snth5RPso7hmfF1fs3axTf4i
I0o4JGMXN8R6m7enrureVdBpe3HEKKZba5Gzt87Igdm7Oa8+Tb6LxLh+ZiRHvFToTBuJd3nDEnbk
MMsZejO3L7zkcnkRM+2VxUksMVzgW4A3bqZ1YBOCbycTziONwpdEADs9LrssTIg11puWl2ZNk8IM
s9E45fN2Gp00939NB0K9JAMXpm8y568yi0zCBmRLR+/KIfHoYEM11RV5KAFMPAvENKarnYgJIxQe
H1gB/wVF2RNwff7hBwZugboA/lTsNxnWVd04eGMy9rRMH746sKdShP2Bi+GFtkeIEhyga9x+h/VI
gh1unQcXEHJloiPyijpAkHcj90y1HUEmOFx0xmtC/p8h4K+ggM0hF+WmGaEWpYJiIIvpuNpJWKWd
XvPWPZTZiqWCuRMgBnqSkOh0fZUVfdPcKROsxiEpbB43+UGXTA8sV5hKtvCtFNtq+OBX7eJgrR9D
ZWBUfCrU5bgm8e7y3GC3SLi5l0LyPManiIMpq4TBkNgr5pVo7qte9Lqlnlz+ys8mcFi8J3qNdgS+
Nk52+0Va8hvItUhLklXGH98RLXAwp2G+LoURgZPkPH71l5rPasWzvjo0V93PhoQQpkuCx7Z5aDer
WLGzq1B2nCT3I3557ES+ZKBTDebLBH9CDEHHNhOrwNHIrgckyftbUXgAfeeq3BQWdQX/RgX0msgS
iIYN4r9HfzPBY7IatB1CM5xjbLJ3zOvd4L2dLO7wkVMEWF5MW5+OHrcsSZGCO8BOdqSvAlQBZyvg
9gebCvU3Pt/CgO2mZwzY5IMESHtsYtbi4bKQPdQlo5bf3zkQgox0SuYrjzZeHB8LOS6CUgl6M/6C
ApNHk0yx64eOu82ixjMsBj77Wzqyk+vkFtgKGi3W/hsqkNp79zT2+FleRHpMF010U9t5rML0FX3n
cHzaByIWi7ivFQpKMUdbkbRnGGBGPh7Drj/eotjIlA/p9/V8XA7Ss3UUCVqvGEh65jeWy9cAR3yx
2I6cbH2vPD+ldRiAzPPXWsarjDwx+zW9quarto1lQBCrZPMKFDKOidFbIGkQ9cMvt8BxdTNBoe6p
Llus5FHPQLl/Ly8NP8qS3XVyiaytB9mcPQZvcpZoGDN95yIexacDZsfIxDEYXpa6Z6yzPt3QR5tU
VhMa8SHzcassooY6ylFT27mybe+4rXdkZoTatBvd/crnfrCQA5YHLgV2CdZypjVcAYPbZsBqkqAG
N8eNewNqcpXJTazIwIsHQ5Z5AcMW6ylQhxVq7X1V2NyqCw4eprcCECuijIZ3HOVF2K441s7Bq2P/
bJ/+Ng05UIdItEzzVT8OOeTQStIT+M5VFYwgxXTMtQ5oG94Kn3QeQG2bkUU0+EYxx0g0nlJLkTpw
24XaAexolb6XnZsVU+cRGyS+RofFTK/hCerL6G7ECAVcs54/INIY9SYNdW2UuLhl6Np3RTREGUly
TyoPTldwkjSwhfQtkPoH/8aqDhVx1DLggBxgDivALQHHY0dFSThi4Goy6QdqdTrDxA7mRGqtYST6
RXaE1H3OmGzjHvX537hvt0B9aijxcfbHqmJ6A38RdahIhPBuEWAhMgdZ1d2tfRQpIppql6cyTQxe
lwfU6Rj8RurHODck4nCEO3pY85Wq+dUF3SuRyN0A2Igwz5f+IOdGi50iYGEXumHcu1oQMmI4xXCB
Xv+rg4QUH5HUKDx/MGKOjIMDahYyBlCaH2UrLv9UtXbh9N1UOWFAvj9zMl1jgSh9o4OBL5E92LLt
7+5pfK4QV4/t7jYduUi4GMM8ibwvwWCH2CTi+AtboKy12H8M3hdQbpj6yQdR8Ox1jRzipYAQe175
6czOA8tcq2FsuZD1L7lfUzECAL95wTDmT0KuqEnMCGPuGSaKbdS8FqX+WJcWRJ/Y5uKxZCx9C72A
+qqe/cBo3S6XahmyY+inoGPPUOliw8cce/ZKHxjOiUU97aWY0VM5eYLVzQtLSfisuP29noPGpweC
9SrEx4jPZhhOqhBOdarXAac7iav+NkQMci3iZJbksrHVqMP7+afkaEJr9Y9CDv3aX5CUnyeYHCxt
gGDu7tmQA5bYi3AcXggjkEvknPeHlgWm9oHQyhJE34Pste6inzSAV1UwMWDWgS2Pw16Xrd4yDW/T
KbOIGvh4AGez/SFVhIlGycscvxLoSWy5ugQlwXUNYqnGA59StGbqHT9DHXrN6LhjMZzUCqSUEZuS
mwdCF2T2Ol7bWD43+sLRuE2eL+jEUaumu6d7Uu2txZRCKjNl2fG9ay49gza2EXpZlVTHJpQCmXZn
ehwp1jA9HQcImZgtOPXLIj8EBt/LA7HeCGSbVKMKjd6ck1P8IiOPhUbEzDHatQFt1xGh5c2ATb4+
eVqhgqcmoifaT1cZx8Gd6sX5utROgH250AJkw3Lh1rq10kzuZzBYGz6W1/7OQEpFHRa5crxWvM8L
0GDaGVv9g6/T3wQX/dHrh+bwbVd6ZYkOp7SQziaizjalKdi2qXabNBY3+XR7XkhrLzeo/FWGZbed
3ln7ZHlOFomK/5pTo26Kvf0wzVA1u42ICgh+XuiV9bC4UyPOsmb7gfXmNrwN9b3GzxlIW0oEuqpH
X1RAnwNWJomrCo4HpxfNodp3uWeHDfTGOz3Sf8ffJw7ncLjaEMrZN1jcsLCei8hq1FzArQdzdxqy
wOI8Jmsc0Nq6nO4JBT1RnxDitwsD9f0dGX4sX/TJussuLehx0DmFsrFx1WvH/3z4+nloB36MRAGT
ZO9u+FIMaUBVKk+aR2LH8SyOVYczVH4X+FsYmTWjkhh4goTqlq+k4dfiWWFrmR1Y0HTpqUiUQE7O
9iOcVTpdVzXk0Fv+7JZzQpTGc7awjTeS1COuVke2P3lXbX4VRoNL+uB1pu++gXaCC4XjRJXtqIRM
OxH7xG9PxCabpAqfiJ5TxVowC0BQOxqTiFndO/JH6kEXYofCSH7kX9bEaysyS6ufJhRofPTPJVJ4
DP4r5FTFWBUY9Nvfilyo6G7vElpcQlhbcWXzerbFGUcEizAnw6boQS7YtW1Stoqo7Hk2cyRBhTBj
YdEo2CB6vKUE4xgQ81MXvQ809bqCh608U7IJU0Ocv1jM+0rLcyViSHnPVSvitunPgK4ELar3wxA/
KO3Yube/WIiBKU38EcA5dCYuCDPl/Cd+9nKtyjUZ9io7uB7JyewhNuDu56cOfznRPL7GNrB4fb4S
PBYWe94JySTNQ/lySAukMckft9EEnI1uuR8DWcAGl1XRIc0MgNA55zRTdeuM441FqFCz7Iyg5XEy
m9c3+SYaBALimIPfxohHV8+s03Wmwm0x+qbX1vIO7HS1o+G+TU4oTCgL/R5S7UE1GUwthTu+dj/O
bCDT0S60Za5qITkdd0kgQq2olg1lklocb4bm/w3bINnSmjqWU1TNktccH7gXz8ap6bCvGIizJMCI
lccFPbpPwaIXru8GFO3kvBexqt6iFpP3Our+MYZmPcaYSRMqjYfTCP0L3a/0mlZUHYhBviK4/vaP
oW6m8Ezj/IMk28SZ+ckBhX06+s9tOr2dzq6m6yhp02YF5yUtjf/oKLD/AYt3jXyoWjOVJTHYaSKv
zzRum9atW4nD2XUgbReVEkCz8Sp2SP6OPTjIFX2FjF8DuguFjp8cdFwUnWOREDXRIyRB8GTICRkd
S/EBMtLj7IupBHxpRbGxduxOsSZOhLEN94RAtLAlbbS+Ep69oPmtA/Luc8OTohPhoOb809hN0/mg
4L2riB7dW9wmJ4ZRI/btZkZwKG5EWLm7SYzl1NIeAmSMFP+Bk3fzxxRoGSNU6Jp0Aiq7PG/U5Dhg
8YUlsqAaOjjzIE/x1jyG324XNBSkUE3moqfTYzGK5H0PuE4sIiXLlZ5igWi+E07i9i4kd3P1SqOz
GWytuE1CG15SGayxEq9NcS3RJVB8Bey8tBHsTpoMiDpPftw1FxoL9HPsUhIkv1qu8nF+2SPriDDt
SWp7J27optOg7OkaRJB6wVUJzstRMt5rxpWl/TPTXWccJGtyxpydZUK0cDnmDAH6T5GTfZg/Xzhr
sPWMJKYOVeAKRED6rsXHCA9IR0CB/99sa4VPfQ2B6BwZuD0yOY7w8+dyMmdF/59v+XhaiW/2J6au
WVelqdHE+EfvQaxhDjb+8lim5d8qoUAH/S3AnrdetAfqoDSvxtxN7lL6hJevZOoV59VQw1LOeLXQ
zgbCR+V7J7WWEE2VRzPQ+Y0RlzW58x5tBv8HivI92LWqHFJ7VwcfHIAtITT+E6ZiNMSrpDH/nlA3
EQfjx+vveYoWcNDylPPVosd2f4K3LcA6MG0jK8U/Rt1BrCkBb4Xcg2f4iyr+ihoRfB/osjw8XqMU
d4EUUYXPWoKu8ecGbHjFOPYrw1j9aYvFyWRcC2+oJPErrvvW4uSXNV0hAr8oMN+Dt5rnESEa/eQi
AlASEHIujtHKA89zozDj8JbywSynpWCBdStcJjznv/c/INEfUcDMKkiPTvMoyVdSNLae9woYGUMU
GE2aPJl3b1M2yMe1bU8rcZm4YP0URljbv6SGe3lKwwu2lGlgf5itILeM383TlU7sfWI38dujXFbt
qKC8O/bNeycFGZszirp+246lY2M3AYgAYGLIhiA3guTx4IdXCxpVySAnKPx7Eju21dKcHySt0gFa
cuycJ6A/EDIjB0ppgRwNfb7tns4vp3+qbWg0aDaBH7yBWhhLSUrs2ezkF6XTPcojnkQkU03hzEap
Aee1JvQrLmEpr9VWM5TWpKulUbEu8/Nadx/vGfDoMTr7C3Vt/0nNAgLFTQsSYMiflJ2idPOjBtpM
bEZPalOrLGDwErIdrh2egX49u97RMnFsFmokbaJchJ3IKGkv+MkziP4UrzSiZKRvymSz+1jp/yPj
rx0a/vq+g6PYc/rXiwmtEgM8kOf3arQTOb6omZWAm2v+EQcNWvBh29TsY7H+izw257iYI/OPrtDJ
qVj5dUEemhz8UKVaCx4JUofObKr7oO6o5pXj/JLszB+iTlA8iNS/b4+4FeH3oLBQIXuxlvQqTpk/
lo/t+hJhYkkIVh54E1C+7agjIrTA58HxlRrQgBspUojz6w23adbc/H9LBrk22ShkJESGl5mZHDv8
mbZ9Alxv2sihsTEstifoEoACsz1dVVv1/YSAaesaBuMLfgzAUsSFcWQnCHui+J9eCVSFSm9G5nb1
YQ2WpIPb0Zxmw5xqH0QnDh6ZYlcI+0h1bOw16/d/01sEU0vmrUBpYv/SRcZCtg1ny2CU5N0N2AGt
8wb17W8+y6V09zMeWF5TjLUq+NesyfytRSRBpElswv3mAXnoqHF6GwWQJzJLQfdfaeHtyvds/sUE
IVeblBKFtklO0103NeT9A8BEPB0DuiQn1TM+zMDkLLMgY3AOyVsrgJeYsDzYBE5fNkxL9a+G2pCI
5bipjEDT7WsomHX6GVr9d8Rr6LLmG6SJ7DxA8rgLysrUmYVhQ+YUYoLPZS64P0mD6TyfSf8e3v+L
1m+g+VmW/7T5kR4JoIkw6sm+R71IOuhli5xy6RTYqx7BPH9ysg6pQ1HUsMx0NLM65YxeDrdAv9jW
j13/Qvvqo6tuj287gvtp76g3fCgFk8psJIwN8L30mfyAkEMez6WYbspAgMFTD8rOLgODQpqqRh8p
6z8VvZzN+yIEbhzvj71Tt2kshO4CiycPo9vSaLYK5GoOnh0y90avGpTpTpb0oWYQwauPkEQzSHe9
dwyUVehmF6XyvtNxmPxrLd2kNytqZ0zqsZ7e7k3+e8Q9cFdcYd2srKR58raI68uFZb71U3Qd4/GY
qr3QhHWASR+xJWXpsxXhwNbd9G1SbQpQ5xeeC2bLY9zMDERzJa1wNLjKIj2UBpiPqQPZ43V5L70j
+Qcijbr/mLfnsu/01EtUqQHWtV+zZ5e8k1pmoae2JC2rmOSlyjWC7OqX3Ma8yiWjarWAOFtNCInQ
UEtdZRTu9Fn/efc4/kTDOqqRFnBL4Oh87nt7Z7/LxZwHiorpo54FJWYlBbv49BDp22jMDPGvT4C3
o2VA8y/GZAcgPKHhskQlEYNQflz9BWBRh8TAO635uAOAEOP3SdbVbZwrVI0cpx3TUprK2gCJXzeL
NSxw1eKhwuIDfZn6nIbUrWLzkmnea0+xZkY0mrGiEokwujqwywyj81qaJIUM4l6w3C2jE2OA0msb
JXXK8nCdGKQ8OsTfMuPsasYXuOF1XJh5JYMNgb+MHLC2Qv1HvmCApFsfD9ixFEa+8U6lSuGILpqU
ueY6vKh8VDh/G/hLSbhHRuZBjoEbMelOlpQQ+Xz1qk4X0eVqp8cQPrldGuSZVjHm69w+5xAYL5uW
o0RlbTjXwr9MQHu0W/5y7GNIVBQxKNUf5GXqze2Pq+/bQ4rlVTVoSbI+nGR71fdY00OLLvwiWZfF
gwXnmmqrrXMMPGu07NCAoKiBd6FXCmWHSqRqlGwcJGgfBiKS08o4w0EvQy5s5jvKSqxI21zLGfuk
LqygMGQrO2H1zxbROIJEggC3PHzt2d8Qv5igM4gbm6fq3Mirw9JIFEGWKf3o8D8H20esvQzg2F+r
uGGNYV3rlSqZdnpNFIsReIJbQm5DW8G4RbGR7aKJ9hYaKGFHRrrkRDameDbx8RrrsEXCyu5/Bcue
uHN/ZyvWhIdWCPoVeu4KqS/bUWlOL9us7zls74s3czM+cLs1EDtmCvqbHMytS+A2wK0fYwS7/neW
Yt+O1xJ7TFdjuHrlqkDuG5qXEEw6WHaDslEXgPvj485jPZtZ0ImMniFh1Np4bEkq3zK3rMXCuDDe
rHTkfkijptW3L7VBVA70QV0JRMIcoJCyNAHEtusCyGTVEYMXoouI5x009kFjNd5QSqSp2HomCn5I
DNbSxQeSw6h/zeIR5gDvNkMZ2tx4mBSeoRyUjy2en2wa3mJIu8SrVnZaOO4qEipTDz0vJbKgXhZC
OFdxfbkGliM2JjXSljEPNUSIUuGe+jJg4L8wDkVAaIp/kDJgOUEw2UMkJjSe+HvmioOSh1ssE0FJ
7iDa/LDADbooEmeCpnZrX+W7i9qih3zznJrdVRriGKlLlB29+Aq6YMqRGh77DzohsbOYZFlSOzV6
55yyxvRbSPvbnSm4VVlqXSmeD9srXFhCTIQf8HwTAe1SEh6P8BEyevhCSRUoSp89fjoL8T3tBtzU
wr2wHxHHlfCBbzjsOLcQKc8hstPfgenXWnF5oPwBEtyvZEvaZgb2FIMFk7T2YswdeVxoaEEn/iih
VZpQTRQyaWuGCHXv5+VzI1tDs49WMS9jvPfawCq4tl0fWBbGGwIKJOaQCEb5a7PfIcfCzPuY8wBD
r/MY7WF/iEsandkQLmdbZIQMKwO/6XqbHE0aMPnQfqcTajzPlsljMS2uLXqeoDOm5KI1KeNYnvN4
a/Dh92rmmke13Wt26eXIVk1fvFz3wDWw31LulU5jw58WBWq5pNXbbL4H/uTwslWe0tG/toH/SGj/
FO5krZKJx02a3WYe7seb5Hq6HkTkLrmS+8/nYSG7OdvFHqXKP46QNmSezzxDQ6f1YMBG7pfJ17Au
mgw9GWcv4e5r2AXdM6FTBw306Kf+nFcTb5aqYbKqQLGh5NQLOBphDWmTGv9I/ZJqJbaCoGfOymWr
yOsB4XAc2CfsMpBO7lus7i4rr5Vg0K2CtnM759xpnJpiDO6O7K0wgl+uufyCpqNuH7a9rpWHpYfc
XlI5jJHip7AofIoTjh6zDuCSZdiXlmwdyjxVEgx6v4p93ooHQkFb6pzJNhFI2WCYCbnw0Lxya0WT
5IHbPx7vZxrqJdz7UgDLsIjClfmyf0VxkY7Q5VO1wRRutuYB01+VPK6w6bItM7lGLnCoYyelkvDy
5Ms6ZAPcSt+dyIgZfjYvvqIgw5ciJ2lPQ8O2gpyffKYtyfl2dF9J0UKp2Ck/7Hhtmi+TxmXanjxs
mgRK3utE8llcsXpB1/CmC2A5itr6FvLIvz39UmRxbrgxiJRiH5HA1r1OiwFTmHSTR70jumJl8EC6
I4un6eWuRHadWgexSfx+0ZYZG6+mWtJymGcTNbLQk+rv2whdRYpG512xthvcJx4czPywYMZqWnjJ
/E71ctmjWM6+HbqVhC9G3jntZFXjm6Md1a5tYqHDTmFKABStfNsyWZP7Q9c/t3YXmjQleongpPlQ
QHciwie9rQBkJFGOZbPl4uqY34G2qRxcIc3u87VU+AueIGe0SSrEawSl3B+QCL28sKK+cA9T1v1K
BcOGBhcH/0BUGNW1ogLPVVIplZGnQhyRTaymXX2RX5u/uyzffjoESZ/8a+nK7G6eO7EHr0x6p8T4
PTo5R5I89uJnE7tK2CR+m66n/qRBpt5Oj4aOmirWb3iC74+QzOa6d99yDvkbZMk4gAV0OyAODOgu
QNrtWCVbqfmkNKZpyVQFbX9yuVp9fY8s+EihgBHIZq5x/IIMER7lI+PKxqoPY3w4YDNUqEzifzNo
ksIjU6+I+AdKsFDUDjb4fED/aDehpsSaCSa19gQObAkI9Ax7iW40FHYsldnjOc4kEhaJY2uVt9vR
ctWoJe8lMYA6sJFmA6MzQZ8PmOnbiT23+dC3NaGzYfcvzq0l2CbS2A5JAOyWFhqYeynV3OQ8euc1
UIxajSXprEoGKpYG4zCg8rl+qJUtIOV3YS9GufVvJQMX85nVa+OUN71l0pjIY8y4p5MTbWobVd4k
giydgpqU+5TcmkTbdWYHYv9CbBOi5USnj+YIyLI2TFzhAL3sdTsW8bl3GTkWiRnnl9Xm4+xkJMc4
Mi8SeFgqoK6c6fCmDSax2UIuLHMYZH+hgQtV54Yqw0YqfKp3hleFqWqiL9D20t0F39FBevOzENiC
WbTmrwZJFVQKxAxsuhHHFxrskLjAYoqi4H01BmN+qexzoZHg+6llE0iWgavZDaiYWVjp0/U22jq+
BDkbWb42osvv/zLdz1jv9YL+hvSslkTAfKWmfNqWPAjw/ly/sx4YtpuL3mrKV7f/cCZB/OJMen7e
lHgG6cpO7oKzCkktlsPznrAeNdEWrIGDdq8M6fImD2LtkOOhJFPCMUHdPSEAiYkkdZsUVO8lDVp/
vabi9XsC48fVd1LV/tFkhjl6gBu0Ya1fFni40W/ZpoyNwoFzy14Z4eYL+UErCz5vYxeS3ntEYrRJ
a+ZuYCpN73FttgcB1n0FC4Th/YRNTWKbvR3kXLMI4v/PWSIvmjKUtBjEqFrCox0ByRNHiRiPLnMY
cwtwzQ1cwGZnRDgSO2zccxwSqEQIEGNSWnGjYVB1co7tWWTwKQqSTBhxLNWwFGAyJtFllCgcJesV
a9AuPdvfAkIHhhF1ZuEsN4lH43Tm0kc8jwSPDcLHLbxaAc/CuOCHIeyU0i0bstWOe/5grP75Z2IH
hg0qloZA+SXK/m8RgiUapfomA+yr3PtEt/Devy3+xDBKRsCMlS+0fslVuXak4TzMQs/lBcVHRUip
xuBGb0/zBDN9f3DUZDNUsGloPPR9/qwc0eXuJm3LTGCJpax9ltzsy3bVdWqvqpvmp5MaqTjM0Zjm
HMrEbCznuGxvrUpWugMZP7nS7bfOR4FtIGGyRM2PHBAHYEfdDtoJ3ajTgO0y+9StHJmeiQ8qHwR0
jA44YSVlJQCxOfaZBP7cgiipm7c0UliuCHwvOefo8JV5pmQyDYTFQPgp1E9zQ8y/ZOtTNfL0DWaD
/eGHPQ6O8cVNfHV0Fq4sJGGwELgDvZKPyXYwwjBHl2kWdVmt9Rc0eY5cLLm7mRgxUh9ZewdBrXM1
Wm3AzCph09zNO5wshDsvTxr1O8yNxyHSxW9VDNraSddCcCPETPS4QNq4XZE3wfaTRhad6rzUxQ7c
8lfiROoIYvaGAX8qWe6+/mWzd5jafzET6l3nvVsUylJPJl7osjbMdquY5EdsT9TsTVbNnfn5Ch5c
5fygsy5cltaa0B+QqDgv2fYuso5Fq99A62dP7Na15ZsJNJ4rgFS/TA8+gidtFRG/cwG1Iw8Tu9WT
r0UQTcjqKFBpxrnghf23GeWixUQyPn9cRvsgP8GbsmduiM3cBANaU3/Vrho7dqvW65vQJBE7+kzb
Hv7ryzvsXKo+9z9EMFDCSuOITRjkYZaJ1Tj/pPQSbhpI5yar8SdNzEURsY75s45O/oi5P5Ytj3sC
isAyek9W9ym+Blr1bMC51+LTs3q33FGQWNECSClMJUzBfsb1n4e8z4qL51GRz+ttOB9yTkKJSmio
MHKB7fJfCUQHlYtT/nEBQsu5LwchUiwR/sOzEk0ivmXh+U12b7Lfuw1yAaj4DUa1/2/swxzMnWYz
JN4pUFgfyf6HaHdFJWF6Rz9sdfxmKzG1XXG4gGRJaxrl90ytLr3rT2FpX10WJ/W1zd6fi9IFWztY
8Gy1CCoegmQDQi4E1wTn6Xhn2oPpR9eXxGjYd5NqJ8N9xeZWBbLgaVA99/eDqNaJ3CvpAQ3Do2et
UY8w3Hp9BEpFAynlvl8oKNi91qqGsc0LlAevsLo0v3DwpiIHxq7SIh/QwXHRGEcMOdJ0yy4Tm5cC
BKul8/r3hiG1Yl5dzkJKs+l4ngqqZETFQzMM44QC8AOrsrriObhG25uK/y43w8yn5nKj/Aj5rnW5
kEYrJy9MbXw7/x8HZfF6y2PvuLzlFZov5E2QkpFkA1ZTCmOE63pQSbFasGg2n6TTE9Llhn4Zbv/A
BafadjT3k6IuF/DnvC1THb4MW+JhQZrsd1bbcQuK5TNI2afTCklDPyIawh5nvc49e27OVC0MMI38
WYcGLNjOlCDfAGs2P9xM4keU1w+ochI3XKI9e8pI+IuQ0Nfvpck6R90nV4xDTNzrPxUzR/zDyBbG
wmWf0pnMYn8eDxuBhQoUBlca2PDpYYhNkiz1AwLbuxA2mZFZdMR6jrow6x6TyHnG94eZo4SbB1Ug
pQxhMHb+pHQJM6ihReDriBnFauuA6S/1hT7uxvTNWn0PYi+zgZcTMJjpmIwg0QRUHlcWf+9qaJVv
VGJI/hz9a6vMvV/WgYxmWYuvn+5YiRFWcta+imNH9wy/xd5SUIbAQcFcx58n9kv0mdGU6zX0PMcm
2aI1a3h+Z6iknXTlIJT9BRq9Ygr+xxh9PHNAf/fFo+EHmpMIA3rXGGfRMVdc6NY8UfwuKAJYj3qn
5wYQwRO2ozpw4Eluxi5sVbAQLZUh22nSW8MYOVnxhVGgHlwjYNwS8m4AGcUgfoLvnIJ8NOiUBD0d
8fjTRISCVPCSToYmfgYG5w5Zn0wRP8aj9ioNfqktIIEiqzJcj54R2j7zALit9xkWNAI9nLxMIWXS
83KrelP5ivICErYYO4fxc+76fR3n65SvILggqJYlB/pifLTc/i5i1RIrEWndTSnOyyRQnOyhmXQt
nGTZ7urjWkUGLpQ7yfBs9RCoHpfVqmFGTglpuitXoLt0Yt35OB1fvhA0VJxYsrWJQFUzYLfZ1NfA
1doMv/2k9IGU8ZSzqhpEbGeRQKcFi3+88blwJWkvr6kALbtOzgUAyvvJfNmtk8lMLLfZIKQ122pD
4MG9gTphBnS+vnrODYgs8d5eUQ84obsD3kraPSpmmlwIVw//z/U4DLzTryNYOT0312Yh6yZTAHEp
hnRoWUS266PQcZpCsAPRfr9R3GitLMT55T+L/m4wVk+YX44Ti/xdTo59gyqbG5sfpBmqZTH897J7
tScxIITbBPS0FnbLSdN8+Z7MjUF72/MrN7Fs8yDsR3L1s8hiTliV2W6YMHDspelv61AUqtaPP+JT
seEmNXDWKTQXftWZYjR6t1xpdpy24REoEsfbIdeP8Wwk6H/cAmyHIOC/7ILubM8EaC9cHTFS/0vi
mzMMufRX/QStsr4x6ctzubIJbpNh/w2LHMRXLc4/r0uc5pMP18pT1NahZiVMFeAdB9o7xyEvtv7l
jgd7jTFESYoBPR6yfs1KLBX7kj544ToQeYPfL+WnSfxyYvwpOotHvoH2nfdjMPuNXGnoDKkQ62e6
wTnHi6rYie83AHvoi/LoEaJZ0LQ2M7SlThokFVSQpBZDibhcpQuKtCndozyl/SlEXL711SzBaZmU
eTPk2Nww3JVkls6m/yqOBtn2NzAg8jsW34QPzdRx3H494Ni0DfbLAba/394skzKQKgznd3tlxXTQ
fCiTpyV6Y153D6wc4dm4jWUaeIlgh38HdNWsmaNhKppOimtOgiwBCtAw9njcP4cgYpS3H8M0y5YW
xp19UeBC4RHqevy+nJYZWDUaRqOAuN8RzNZRJ/5fNdZSyUtsH5sdaoI0hcHppCfeABqPkgXXTTxY
6kNreL6lghEPeQSJCbrZ8OvvNKkO7qqR21UJz3pohppoEZ/iYB1N8DiUIbC/XHykPE/oTsRZlX8Q
pBSRzxO7XTTkwDgU03aQ+ed+8BcOq/yKnny0rcqy2yH1QAoJGC0sWs5+SngeZFjQsVD4utq3hSD/
g4ViGmbnEtk3U2uKnGfkBDj5TdcxHZ3saNBn8l97dnhP2BSi2XodEtAunz/QosV0fhbaOjWkEJb0
dKJAOVjtw853yhK4K2oqtso0YAg4qTBjLtVA/+A/ujC1it/QDio+jsC42IWjoRLFkBiC62/WLl13
C72KUxWm2bZI0GkhWqiETPK67d9sgAHPiW5zL3fQUgVhwFB42X1d+/0maAJYeMv8XZStqMUBIuk5
6pHgI7YVzoclt54bDlIoX9wOI/SuqF7b3xX8Sz2NWfz4L7EUgMiHlz7Byo958d6eo7qJVnERGhjt
qKTBYc52dsfz56m5yXbQuIP6iSYg/4dWq2EhCVPavOB+Z+on6n93sYxRWAnKJ6KRnZ6XsAWZl3Wb
AjSK3j4nz/y6x9dG6/VY+NzuJQNi5b5yOKi0St70HGTzPVGzWKlBCj+Vz1PzUdhlXOzdn0DYA7AH
3LdDlLyMjF6YgfDD1Fc84WJkhQMIsLUq9O/wDIGomoPyquP7UNhKLjI+NJjoRo43WRFDz6XVMxLQ
ck/mnvDraM5zgIrBJtAJuIs3xQ6X+O/Elku3sHb14ze+3UQo2r7tg19MZbAR57TGTpxIcKSZ0Obn
vyJgOLJPif2nACncq36o0fRapwkyN+atcAZqvwTLUSkALeZDh5JixtAtc1Yv/kPpMEJzKX1dZE/b
7cRUgs7DFMNuAeMZvjjr+8M+h3JdR79jHn5KYHZVvtQP5fLZrM89uks5Y0uWrE+gsmX7EN1huYN9
Xk4POcVXhH/h2EO7n8DTRHHL+iBUM+xKP4Sm6zv5KQjyHJcJstRPvL5vpSDLTqJ3zMnMQkkXQTF8
QZaYgfTS3JrkINzN9uaPUZuL+e6e5bI00KfPhzQgLTsOdTiU5R3lzM2AGPpQRlPjeIzjsHphS1YU
G/hUTXcRotDMkvujb9qleNX6lsgUSDmU6sXrdL5eLa6cRdyFIjF1QSR2lA/WVRq036dNZlNuYv5h
jIeU67PUaIuY2ipzCxmQcmBA6pHC/P+hu4skU+mcHCm+iJmsvhyaiU67bEjy6JAuMT/BuzE1L2hT
Awzv1iR+wRoOQYTknsFZC5tapSsTsKj0G5B7kfSCisQ3MgMgTqjhL6J6lo4wtmuy7RXmQh247txo
qZyVgxWpzdrVbRTbhwtM8fsE0fyc2f6u7zbzbWIHOUpRJ/5Roh5ng7HCeYCv+E8jmIE57Le0ktDY
fN+P1Qafw/KK+JpuPYf3M92nURmyz56gNlnmdurYowxxbUywlvdrwIjt4vHM0uC/QWZrKgRgnch+
5h+njxtQObHSb7ye3tPjcQREV9uqwqJQ0phSkVXy+0FyXgStDs9zoyiLuqqjvV9zYE1b1ztD0sKX
vrYZJV2MAiVJG/Sc9AXkB4qEuAaw+P4v16XNpZLyGIwu5XYpWH3Ho6oFzqgLBLDmOgJESYuzGxcs
IihvD3mfzDgrWJxFvbiqQw2EYgS/jT0uKoBxJmQOM4BUOdT+Dw2Hvk0R4KQ8Qg8fGCXkM2Rzf2nt
XZXohYDliRA3J0Nd6122CFIzYl7i+gNceFoPolHorC0usXB7rXJJ+NTl6VBJzN5s1RogabuVc0qm
WZminKJGcWj692HnZdsptI5KL2UnVNdDVhVzsCIU+v6qDsrtyz8UTG18jSiyzoiC58eefu3m27RF
zi2LayAaJi1Neduq8JfktaaAvu/si7ZLx2rnM0j3kRUQAI9jkt5JJ+a1h/85YL3FZ3IOc+1STMut
I23hxIlN7HdG9Jga3uthb8w+rgaYO0PgIMqHsVJyJGLKqBvR8aYZUMEVHNEZVrEWEN+6rAtZBd/T
+n3DkWi3tLSc8+dZG73BGXK9KqhNpoPT4oKTp53+bGAG5dntpFkwvuDLfCYXXZ/xHd0iZp10wGJt
yKPCHh/eI+RtANPLXTfcvPkT4cR5RqzhoR2aQg39LSoWtG4yBvA+uo9VHDTwTzMCXMWDrmBS9Fby
rIqtm6S2Qd9zug5s2O2xyYoZeYO34MdERo516aRFOadG97D955fVoU3duNNaTwl//I/KD4N2chxc
WqSm5w8DMQ/R+uwYHez/NQfeXUy9jR7XjbIyB+NR3l8WG12ElM/uJPst1hzR7F4o4dUNwXnTkPZN
BTT9AfTQYnJiwJQJiA2MMMFRxSAeBgfthMVDK8lPOBG3gpre1843xvCpYqSokssUJ6Mb3gtwX1SS
AbhXP49uqqyCLNMydbmA8oGaMuJI8iL6uva3A2FHDJodS6FLCPS21LpHUb0hfFBugMnCphCFtM74
1X0ASGIrHoTRbYXrgCkwsKq8+JO03OjvpBg1r0svCaJC8BOeWRk/EenJ+47reTBfwTnX/Esi1+4b
CcaBEKPIpUV7QY9ZhF1Vm2Blr1SWXBYTXy2Orgmu9U74sdm2xdLFUkdMlvt0BM3lorDZ+KXun/kx
GaHNgixTfWo0S9I8RSZ6YX1nHvSuTX3hwD3jplFIJdLcA0pA8rOFNFzTANh9/O7rlOpGO/TrF2tx
Hc02LnTRPieXPPVO7DTYQ3OKShtFob115ERYDv9oxd4vVgdC7TQEY7DTtmZEl3dxt+KdRCJS62cb
zKcNfQ+RMkuZ3vstzIjkSq7Kzrqq5YvOWwpwG1b22u1zD5AwKGmDEIT5OsZGJo5kbSOrowMXNwER
xW2+c+1fnjF7UKXfwOaNcKsCtUeWkyOdbUM5f2lgb6vkNRxOBjr9nme889up02i1gyp1cmUnve94
lW6QhylFtDJI263s3C+121xb68kdhiaUj+dWZiLpt1cU7O4j8vA/jUjYhqBHc/Ls6ujyUxzrvY4O
L3Q7WaZSC22ZYut/iHolx5tzLkkh3uFuuvnKB3suHpLQO/rHgA1Pe2mGihUhseJjkiGLpQAxQmuG
OWBz75JX3Lsv4VXQEM45A1868JlhrJ1qSWScjYIa9He7uFvPM580fnPpGLigxP4qr2GzrjkhK4M+
fzV5JzNPF9mRbYISLnHb6brXHpWg66/lAFKXJydi3F+3GAJvCbP4NWUIUD5NFdT/lWQxojO0jOlI
ojUgs27x4JbG2xUCbo/DAtihkDQseEtxR4A+kwCME/oFmh2U8iniR8rT/mzWMGeNn+cuZYT+r61Q
yoh/0QZHyQbigrac/cGWfg7bsS+tAhwHjJlK9zLVbVTICoNXSjcqUDvvSZJKuxU/5wmCXKCI8atI
ix03VxwY9oQtyGRU8NrgfqKIaB2UWVGBLCry6Q7Qk6LKEmaASQYmiOppnxzTBz2vuX99Rt3OLYws
uFfMZMyYzJ7UPYc+CGtBtgjUc+vHnkxlT1iTfYbTuqE7QMPLSAh8DAMUOVfJ0mBEAQNu5a8bJ3vM
CHo04f3DEOorqOn09YnIYrtmbvkjU/0qkkZF2YxIJCLQTrI7Sugq8wVp9FXEzuKKwnTWNh4KCSOR
UfCPA7uvPLxuBHsmZ7RIrn3fdW4Wyd+a8tIHdb378LWpEVwnL7va2afWYDj7B++gcj+pg1sUnh1Q
kR+6UlnDfAtqndQQhO1Q4cAwTd8N0zDHejnFpSS+uyiaU8eZE1NsePH6ICIQqBbuTngBVdwjaJKC
rGSl2OHzmGckkreL3jthexpZwWzWvAZ/jVa0qNblQSUNSNtYuULwaPphAeD34BJ7FNNz/QFSaAMD
Au4JVdCPRK5lyPtDiNVQq/fPu2G2DjJYx/bi6OtPCHRVLTpdjUuOSll2FUdIyKloeCOqJWKLFuHt
4eEB/jFMROjA7mJ4R7Du8mHWU2ZgmDBdo2gYZ0468YwhSDQ0pzhJaXPNTMsiO8RHFWXLDoQ0bLrg
Jh3DBIsVsCIl6nxtut4tgmo3YJJ/re2BKlKOQwjX5bwJLrrk7EvU2eIdclQO+AqkZVb2iPzXPNh4
1wD68MDgIUFxM8ENvF/pg8EGsFmL3NHcHIyEs3vdr6xSDCdZhE4jeOOJRRzIKmkh+iAoTNKwzs6v
IJlcpCPCg9Tt+MfvZWp2/wS3GmfrWTbdsGRdOJqOVRFNkM+hIU6CofzioH4TGKjyOmwPSgJqzFS8
t8CM7xCpV4/8O2xhoD9OD2UNLgvRpWUlnBlMMuTYiC+h2/s0YGu0UbP5tZmXaAVRgqY4aV21o5XM
yn0EeDJS/6O+taOO/PfzOxFWvwXAytSw+tVI8Y8xjfVzvYIyFfzqVtstbmdJBvloI0PSZ0ZIEO+D
dO4jYv3DL82Tgk+QaCuKmyDgiGE225YmneJb1cb2ftaxusgcZVd5IxNuPgf8BJGgCVedxs8maWm1
ptcdsr0bIkq8oRexf0H19yeH03EoHH5bFYb8C4h4kRFQdhangu2YHNEAsG3WV8tkuXzrUv4XpM0U
weicoAPIP0jcU7SJxlZDPY4vyr7c7x6qUm9rYgsJMS+BoPHGDPe6fVNstgVW1AAaiSyoibX0a0DX
HkHh0CIPl0eA5RUAvZFq4d449CxPDRapKwGoo3EmT6hvSN0+8ld1pCp6/GdMBAOmT+eO/upQk+lN
Rdwt++YzQia41MQV/RjQ80R809xNEEuRTcKAdOIP3UkDu1mHY4l5ldD8cEMtW3LH2MJLHPnRWA8r
1DlNKHBjCpbeAcfMyWqO+xdGf9CwyD6fP326l7A+z7cYBNa+oRgO0GbrpBhHqzOx3FfCP3B8wBw7
5H2tqZbne5SrHPplSZdTJ2uSGTirgt0e9YFr9+TnSJAP7Iy75C6cQ3AZjVtIh4wDVJNF3yOzZJp5
eDf6U168bFAjuzfMqhSm3sO5HMtTxCWP+bAjwkOeqlACgR4kpsOw2JbjWzFZjzpKmgU3JVFWgGNG
5uwRTfUhkGs4NJvj5H+266xIGRBWH3IYacRFouc1nRnsS9PXneOkbm5BP4nhL2+w5OWRP6K4OUEo
fqCpNVcVaaHhu1pF1R1zU+ODM+NcTVpOejlCYcmx+Bwx2+A0fss3aPv7n7d5WW9cuAqwXm2W5+Oy
Vp68Wooz9QAaFRyV8/3JUQ9z5TFDi9tLL6Jbz1KSx1rL5t1tyVgPuHHIrMFiz21D1hjCLFVJ6X64
DrcCn6OE4UXdGu01Er8UmlGe+OeuqXyKvayi3w3KrSMK6+xr4ZKA1rxKqZCox+N0nfbqyy5mBmGK
a4rzCpGilfOLjBWpEQcXcAfJ4Dokwv4cnPGouiCZ0aTCxmJx911/CkuekMl7tGDO5NC6iaiEWQYi
VZZJ0hrWepaJT3knGoAnQhSQrYCXc8PvWHnDh/1iSlljSFx/ajY7FtrmOGde/3NOe+99cLqXyT70
TCMMrN18dH7z4WaO6C3+FEKW8LcpSyHhzflHpl28oAhbn13YpcMuep0lsxhVpAUqGPYqbqwh0ihV
+3WkO/AbP6PpbOjYLOmJ+xggtLzB+CNLn/IQNNcpVm1CmIu3Xe/2PssvbC2cnNKVqtUiEbPVzkVY
ew+dV+J8vn6Ck0q9IJeQHlJOGeM/IukVf1N4bq1n8/Jh0r0B+bzdXkzKBaJmH1c43A04kcaI66Ij
SO3DwJmpXxFzSUsPEnMmEuYKmWr2yWGYtCQ1WgE0DN940pBnESr5sCTCjZvsRBMBz4q2uFnLcyho
/dT5ZItQc6TAX+twJ7hoLeWYMaLAWOsAYznt7gHcB0vFmB63mburlTM9d3ASEj2DTJ1rOKDB6Re0
LABpbSYhtw8ZHE5wYTPCZkBKeXX3WzSNJNLJutoxVhLd2SYPCWODsaDS2Xgz7ogqk/yYlxpxSacy
XPcPfN29mNRl/GfQsM8NyfD9vt5Rz/4h/sO2xLxfyItZ4vNLi6hALaq6vZsBDPO5bSkSuknQooYj
IXS3H/5a3rnxcn83J3+/rggVMgeSXPZsXZh+fe/fPdo8m84Ej+n40XiSwQMr2I3X98Pg2T5U/QQV
jXvN2UtFkMb1bj4gbgld4GPfW83n6t2qfBd9BukyHc3ZtB4AdaoAlFERTSmii+3vuwRW7CI9Bwfs
tES9O8i9cvcoGeykjhHfwez5LPTHEGNH/6m7eC6V5CoCH18OeuLlWIDgP3xP+ZwJf5yh7HnK4baN
FDYdweWubcrkr4tyut66IGGNDyolIZ2ucEwwYWvIDBE7yrgzAHCXOkTvVoAgB/KPLIvyWQG9aBrM
95mUfuaTewlGb1rgj6nloj6V8fswg7jtScHetse1iTfW8Pwrwv8dYxi2D3uIp/4FoIe89/svSLHU
XkEHud31KPZi7KoeCQ8vL2UJSewKuSpFbcSdAntbvkKzcKsp4YqlCMAtrqMG6ALTRo4gaYVRt64q
VGwuUxhGvso1BkKSb4vgb8K9vbEU0pZ/4QciPS0I2oijxhaCM0mqA1CHo4vU9ScPBg5vAsAA5qjj
iirBS7eCBSDYxjMXC43TObzFFVMAl0jXD26az95Y6fEdjFssonjWwRDvOUF1MlDszRpzWHMcakAL
TdVNTYquSIwwm4ekhIzLAIy0c4T2/ASBmwbgf2Qxn8yIEi6VAEki5DVdI4XpjVzU/11OnZQ+Z0Da
Q8W1Sqy6wMOQYOqjG09cXWehvl6/6LWeydxZ8mGlD78bKrmznPRFKXucBk7bHKoh+F6HXtVnUHQX
ZI8BVuDgmk95mVOd1Z2ugd9XcfflEVKuTVS9FwMul6Q9KLBTtkfAugoIS//oz91SpjdC89s4IAQe
MwgSxS45BIt6kTGBu13t8BFL2+uWYqvanbvD4iQZqDxHhXig442WcWAuHoYsIMeQwI14z01U0nyz
XndTilLBCDi/G6zr3Is9DktLYaqAzmiuXoIVSUbMARg6zdKVvWIQn/Wp3uGPjei41PTIspD4n7eZ
lMREjkAHlNk0CzrModQfbG/plE2WLnPE5JFv7gmPSLKyNyUqttP12zDFgHJ1Cjjw7H5iwwCF1RI5
zxNemTlQotb0SWp20De3U/Qs5rOj8WxicO++1FNxqjWPgJT9s/RXpd0RvzLS1Oj4ZOI6w3Nu3b/I
7izJOAW4rcLra7ZFMc5drxUp3EfnpBT2lwKokOLbJfcWV5iwZyVCKIkuZjv0T+N75Cwd8t0QWO7Y
m8SfC85hEbtKKn+bZhaIBy3BRZWoiEWXv8NICaib5TkQkD6+5l7tw/YxuajxYxg56Z27yB3Veb6r
x2D38+erouqiG/gy2CaPad04G23PIXmuI1PHXvJlv+UfFt8AiJwH55e+3VRl1SnmKfTDrIhr8S4z
b9jsXdHFJlM5790LWNvBmfIKdCY6vkt/Ej4KfRZa9a7IZfM0VDvFXNNQy1Nb0pwdHnZkoRUIljU5
8/zI0kDLwKJOFcE+d/8cn4RE+lo3gzxP4rbobns5WKEud8m7AWUMlDfMxACuDoAHvhrXZrcHVdNE
SLLkCl+pXvbEL/2z3hfRsepEVXPHaMkIwg6MN70Chi4iRuLb/lhqkuFMHYXdOFugi8kWHZsTFigG
TqOlTJRwEiMBA2btcFTUunbiUZj2RZrCfYsYi8RzFgD3yDjgNw5wLl20NQzjt8e2neRJNe40H3kB
vPo/JTag59Mhifn0qjcM0V/CXiskCL2Jv61c/4ojf+CwYG8oqHc4SNiX3O3M6KppOC0KOfVZtWwi
zhqNhkoEwRQEmSHO+FsACxGyaZwVpa7mAwKa08UU3AHrQz6maHg7zX3SSW4nQ71C3OSQS80lJqCX
h4lMGyHX9XP02KB7wDtVGRMyDA3J5ODIafBC5lZKboBWwhSpzm/jKVQipSCUQsBe3YIWWh9hV3vI
NEhfPNjeP96MzbyR4gLJDPZIaxmjRUqPzKjRblNxM8J9IhY21jJN/zfNGrWWebgg1oJRQxalRiCz
qfJcvM2ggwgJ7KaCX0N8UHHh454gUxNJK9xy2T2ORBUP/rEUYR0LNFBk/9ch2Ae3kmRyzrOQhPF4
PGhVl3tea0i/Lp+RUi22sevYv9bhFxlqGO7UBbkTHOyr0WzLRhvCNUiOW/edlScfOvvBH+atbF8C
Qv6z9uDR1L3W3eJR/+tEXiYuOW8B1nC3+HH+xKnodNDTy1GQMc1JvQod3Hbkg1JfxSNk0RU0WpZ7
a0DNsyg5aJy8pgyIYelJZRg/sOIhAd+C1zaAJIwrFi17xNwNxbKKpxkwK9HoVPc9sbn1bWEVJgaq
xGoSEKBsfJFhmjzBby/uwDBZGs07qj7nmCMCOVzR/lVHyqgF+u9QJwgWvOWB5D3yIfiIQA/sVL9u
7KzXzPssUNsgjkoN9dMx4TnECwoput4e0GIkrqosnzJM0hoyc4MiN4DeXFn+9R9jHzHt05YQpdXu
/tbIGhU8RZYEuYNhnTrhf4efKqCfJVuqMCi+QuQ12gz2B+FZDGZbesudlrw7QGcafcU9dH+pmrea
bYDdidMohmuCYX1OFi2cdN309jLQGCejKXZ7na6MnvHdc7p+iu2/7suk2kCtAF9pq64g/2mdFbbl
PEmX33jXHljQdTmxcgZDEuiq88WjbZoUyTULHfINwLlXkZ7CvalYCJbdHKNAvAAkc4Y6ukeMKY1c
msS/eZZJ1YxuMyP1G850nqpu5/y5e2EpOsxsT0aMA1pgB7GIHE90INCOTprr2kIUmkHRIPqAQ1cf
qaOnMUhjv/kRYf64SsIsSsNvBvI5gkHspwbvTMxNv7lnGvDtYhPHmo18h97EoyQSD981d3MtSikK
bvGKSZ9HdrXLrmyUuJFvG2WlvDyI/SDAjQW+x4PiOki1iIqxk0xX9FpxJo976H+u0iy622C5OStp
xvsEv7sxe67q8L5u/qdGMz/yQ5WRMrMdbSYLpY7Hvj5q2xCGd9l2yU1lELEbvTSceeZ5WTliphSJ
uACoPWu6GO2KQKnI45sacuxuMyUnkk1dbEv2EeHXVRbk1WwmX2to9/S2OuSJ/D7RrQu7GwUbS7WL
WhRCYjmRShiHoOpsdAPKt4GZh2/GOHJ+nHDe1y+le7Z3mF7L5Hf0k/nphygcA13qbU4OrieiPx7i
QQcu+H4qMGLvYVIFFCl/dqTebjDieC5HXGPZRfp7c/LqpSxn3a5U0A+F8Qp02L8nz2DnAKOASffx
dW2f2m+h0d7uLkBXYGGD4J8gpLMIZWcTYpS6qIMIW/NCK96Kp1M8YSIMDII9NjS+lZcB50DgoHXt
r0h8e6ZTZ+e+diUFTaJSXzjmpbojEQr5RaQ51sRWLIXLtwNR0d5uPfPGq+OZaKOsof9Z9n3JtfxX
OVrv8DMq9C2KWG/V7ICCTHIUZiqZnAklmTxHiFXv1mmZbAhPpbUzyXdpnFrlOHSDP0cbHFlP2L+1
g5Bhmk3FM+OGyCDjUob4/Unu7gtQRqxWA2/pmr6NRNybE0j8n/RCIZkNCf+gjAtyJTcPQYV/jpfP
4qLs157pcdZvuSWqfwY2JxtOFDRB+fI42ROivT6sR1upemKfTdUnfkG7vu/cxpJlcRs//C2ETsE5
JxjS1suz8KDWlpI5lXuBDTaznPSRgnBCy+sRx6IZ6/GK3NsmdTiNJNxzab2ZUfXyqEgkRRswy1Y4
cxOqvfNidCbCPmZO41NjcFl8e+YFeqngueSizyyBSu5hw/ZLe3VChpIOA5+Tl+Eid9g7zjLjEpw/
tS+IWT5xbOzELn9c9vuGfiOgiVCnfrA2LwJEYeR/itLzKQy9XbkSBcBXmRD8uynr6iI/77O5Oo65
EWGyGAWXcV34Vg3yHz8gzm4MBwpfQow2Q0qauV/k+drNQZI1ye6ar/br4drGzOmOfMzv04J2aC3E
FffL7MerhToB5g4qeMJvLbkZZudHyIHmpJ1MWTsqjxjvkGhc0qx1orr0mwYBEudSpYELFkDFrVsd
8ddvFj5UqHBykJKdUXL/ureiciIWgloAaRkjwX0CuWllvw9Vcvpv/JMdCnjIBHKXWVw3BuVZWN2Q
hnYV0uaaDXywC1Rxpw9Rc6T/h4c6EDivvLySv+jrKAqHuuWTqw8h5D8xsikigbeVkq/YU15JSgE1
lue0PfD8ZIa8H2Ohuoi503iyPemj+BpLS75aH0p3/388MDyZ3GJbo3QO1XXeX+qawQ7KTU1Z8VqC
gbnZcx4oprLjiTKoyNOYWMAH7mf+b4Bda9iiCZa8K23UCmFkDWcRlvo1+qhkSaFrCMlQTdLf3Eb6
BJGWeO3kzY8v1mo8V/BmSmY5VjN4HXXHS0PpTM48GQfsGWzH+DQXlPBgXyySOU0ytcJNLHuie+zj
civ5GA2+19RvPLY4sVVeTPOCzqBoEEdZ8uByBIvRAaAkbULfEulg0Y3i0MPsTic9xcgbicjwadU+
LESgkgf/oJ1GGMyUo9rZxo/lRGmT+ruSwdX9/619LZwVYFSpFbXK1+QIvySFbXXbYJFshbWHFkeh
WhXg5TplXYIuptmNYuDKyLAY8YqUkbF5ZiTH6eRXAW24bRzudZNQsq7+pPcEJUp1SEiNWgSmWrk1
1TpeT2gwso21eT1Kw4UZNfoquuaSexRxpyf8/FqiiMV2d5A3jyJaXzDl31jzWT4W+yjwKumdWsMU
AOLAIvmiivmdXaUfzTJYhZieCgUdRjcK/mfPD7mA6VX2lwC37l42hq1tvslXi7Z6j3xs5b+//Nfg
1O1p0D1CKK+JB1MSvmIM/09Pd1589bJhxOQ5cXZBmJ/09CnPXmDB6Cv4oMKMLpJVxqnyir6zq72g
cx12a836YdSkZ35VFKMJYWz5MdPLNE4HGzy0tIbDTW+CagvgCKYv0alfQ6cUcutdPW4z+62AJ0mK
i/dySXCpeQTO211QrVG1EdFVqb2o6em4wF3/29D17CDQNomUtrZq2/B4j+MXjkq97oajKpHQh42z
djoXIlv54HcKGTcs6/wtalSaHbaJjhzz+eXL/eX3HW4hKOjiNtVBxCpbtvejZRNORKVDsY92GaHx
ZgQ/w3gzV7ft1frVIkL+q3wx09KkPeM5w5pmi2Yvo8Q1ZeFYYsBUtwuU9jJisyBj3RB8yx2436M2
K3+2UYltcU9pcnwmVUDtVlFDGtHe6UiVjgJEPsSgYPydjsiFtc+ynE5NYzIosjzg3z/thKFA5UG1
zD6O8CAZT4tkSMnSiel9u/I9pVja4IkIx8dbHVE2kXh0LcYprPOAg4/NWOqngNonfJPyJxj3Fwvt
bBdXJu42h+Ve81PoSH+izbkMczIkCm56FMOl4zpE6E8N4CraMJjDtVSO5GpdN8u2eTw2yuhxXQtP
X67l/s/VtMyj5W0iWzx3pEyV2idCSGjXdgqNFM1me78UDJazUjYjPp9DKVSkEKAizmh5+mO/Pyye
/bfHM+0aCF15ItC3+btWYFMbPtnEoWFCdPd4I0DNU4FX/ewsNTA5b1qMINDPqbWhneCQUXC9hYJw
Aq6pQcH1lp69pd7SBJIh9nL0grteggNDw/ErlD0UewwpD8CIRIAjmP4qf3xeAGY2w0xlNR6AMUVy
SNMfRfqhxXWl2AoTqcHtAF0/Ad9T43udvv2dXY73n6aauZQBDPxtu4DF6ZKH3RqK4FjafbE1wAPj
CEqu494j5Hnid5ZOYVvtXbZffAU2opLDbAq1b4wI61uO3f4IIMeS+Am+K2UDDSlJiGGsj3YTQAXD
PPNQWY7FyA1uFFCBV8M6MtUF7h/2LpUzd7iY7anUJYfIiFdW/t/DEBl+DaZDrDG5ii+ICOO5gJFg
HAjqAU8iUfpzuLdv10ryr6ensKl1tjoq70Nadb6RTDPmXt/PnxxZZZ1jNQuFQDoGXdiTZ3k6GYm5
Zm/VJcqKpSXWxOfVdtKydqBY8c8yLhSQZ42Uu0sRbiXcQNp8bgD28l4Rto/IY6bggy75VkiyVqHI
rcjfKL8DRDvdzOCNKVHRB2JHNwtrXhMZUI4FG0nKLKCZdvAMLmxLKVsG90F5CiZexdw6ce5uEPwe
0y0Dc7RXAo0G779/dD076tlTAAsy+4HBIPHTalrZYR1XwMeKGDcaYF7XOdZ1l8mJkXZdLYRXDVwD
L4zAK7mw/YEmmBw8V9rpwoCNnXm39rCRRZFCUaN/HPVc5PIuMi6K3fHfSL0aWYapmMFSyfT34uL+
2pozIkpPTxMZ/IF+JNI3caMY+yt9Sdve02I8SYUIcr71fzD8mplY/FfDUGqYYpKtaqUa7rzN2jpB
sjPtgUgj1jD4bYY8LtdOG2tPtN3etgrIRZBD/PwyJq82vSiHjp47cQ5ZpGygWdHdJ2CDkRIH4t/L
n4QieEEjbCdufskY+x9+c9y7MEBsq6BxhyKgayUOYVmWHXY8MhAMov6bNDM1nqQhxel/lwXRy189
DTTrehUSs1piB80iRaDjrBHAb7d7H8vjdURv5C+er0ZAnOWZcNUUPwdhHjPcJ7/Q42PQRU/XO7Mj
zV0JmKBdQWEd+VImfe/kABGpqgncgE1fy9ISDeRSITRqskaNKjJio6V2QUapUIBlAzoq1Et+sBY8
CpCu15yZjKBv3YMjI58gCkadlTSMdZCeGD75HtmGSDIzMUTqe0g6HOofihuUojStO9yctPrUViRK
2D9AkMhGuWR+oSYa+QbgvR8ddVVhMpSaxJ8kqL1gbFUDNHwPk8TibVRA99/bUnSc8JAgCk6bnfOQ
sITr7e89zjOjoMyQ8J7CKea8gZytwBkFVHwLR2wmOptRrJvTgrNUezF3/qvKgam4RAlmER13IM5F
ZnAwxTP8xDcFhGPguvkllo1+k0aOuHYRtCSONGkgzmp0IPxsgkTrNjRXsyvxh+DgBzVMzIDolBxl
dmVZoVMdMJbI9KiNBeF9u8D9NnxeJ65GuNxJr/o7ve8a9kC/fORohDJBt0VhBW/y5RJXgluMqO9k
xe42aPJSNq7Iov+/FnrUiKohpJuk/kwh9xlzeBgMoHE8wUfovIxpWT48TgzbwluGykGOvBeBzro7
vceDpFeF1Rkxn73d3zqvMpoxeyGm5nKofPjF0V8fKYWzA3MZK5XvB9WrhckI3Gwn4dHxPkwiGPEx
18Mnh6IM96JRiFMNYMxsPyd47dayG6Qe0t2R7wB0/k6ogPI+Zz9XZej/TiJ4QqaF8aYWUpdzI8lK
BsxWuL2Fwf/H1Tul7ILo1uysASr71eFqjMzv1zD8j5rFBCl8f/UJA3+h3fZRfkUx9odFqn8UCC+I
f7swLfRGMgxfNrfZ39+SrFxnMPpvSC0mfvu5UahD3iZGo5ueOYhscMC/ebeMATRCrQW1jaFe5Wx9
jCvZgIJoNW5XL/i4qmycQVlvyG/jph60OvvZCcKzzrwZ8+gnpjNy61zYp9DUjq6AOWGdc/1AXsGm
2fKqB1L6KEzvZsdL+HBQkj7vPW5KDACqPsriE5BHTR17dPTJzA936uYhLl0SPmXnKk2TpiK5mYEI
u46wpSb11Qjbr2XD985mcCdeSUAF84+DtU+BTE1IQTDLcJHOJt8TohvlFsPiRoeP9luB8M2HDmyZ
+zjEgXANpcqSW6fASO/vlE1cGxZCkLK3PZ86gbHDPXv8rZesQVl3s2GR8OktBM0WQhq1OLr/0dLY
fJwVVRLsil4WbPHiGyi4KnxGxVl4Mw0EauFMLH3RXrEDy+pAvsZ6ddqP2OEsuHVB7btz1B0KzLt6
+4LTWtEDl7SlIRmo27qUWUxMs3Mx5K5WQfsiZuJpQw53/27RxoSsuSroIXNVGhuHi6P/+gTP6fpo
6l1uQozL8qFDm8Weqiblyfm2FKi6Hm8Ph86TB8mgdtQfAupKrOJQMY0X//THZkFarrkBM0+YAP3f
+6dg0ChCuX/2MPQ9/FV8wG/C7jPND3UgCnGMha0QSM+MkVxRv0/y3V0vNDhMWCCm8VBHQesevRa7
U9LJTxhOB19/nJ/kEVKB0And9DehA2KJWVkuCYcBDKUq57kialpteraK/FIiadaU+GhcvxBVX+eg
objlIcFueCWwbQmAJbOeTLE/HFtjvSIeMbTJ40147xIIoZa9WqdiyeX4KoJT8hTrOkhnv8nctDfs
mN+mTEj9POAJJtFqxmFCUhoHlP0phzuWilXNLHDysTXm81Sn/c7YCdZc0A6lFTQFQvyavMI0j13m
nvIFclCHox1wf2YKmhl1YfGq7p9tstEeh4L1bVNoFeyV6RfpWBgf8cnhLAjpbpWkfEwKB8QnTdaH
zyuGwE2PY61bOP/hD/tYBCBz/zyfgFY8V5ngnEoTgsgOUw+hAVzry4wQh1OzO3twB1ors+uPHp2N
bIETTskz9d9xV1KIkY2kmKfQ8sKhu/IMfQZfPHYnzIyRVg5y7FO5n7239DXujS3n9BuqyH9hOLX3
wbY1iGWFQlE0VYy8Y5EzmJtK3pZPe8BQmUspfZYpd7fYXR3b8u8hOkkQI/GNe9vaLJJNnrraL0lN
PnF88vlY5FtFfMKBOaFvdhiZ/IK0LiMeocXFAGK3N1mhXyTZFOmSb/wCx6jk2ZfYAz3bwB6upEy5
KiHT8mXblLV44KwKJDSwpOoidGNwEHT4ZqU7iDBvqt8DMVa3OMrImuROOnsEnUK5QKJotiNxf9IV
FdAsHdAzWtaHLRpBoFwpu9qiIYY0v8RckUeuK1khcCee8acIQu4NtoZpyR3oP5ebEJrzZPkbSAvU
hblxLIKjiAqSqaUCndnvHHApV+cLUHKdbjRPeEcldY1k+AqinQx0Q7oT4+KpwGPISjn4+agjbI/q
5IxPlCGgXgqPuhnV+9qtwtDQWWoT9C38NA1hS1ATAxJEm2H6aejZXC6Y1zfzTpmQ0n/esEEJq9Ep
xQO+MoHPno76LxM8HNuqtvIjWx1jtJrpNt6aPQOdYYqQn08oTB52CqODcP8RuOuS2ahkFnRuZHGO
OkRqZei6qov7Ill4Fo/22qMC9tNmeco85EGmVdUu7cOoWYEKyaSSyNmMr5SlBwWG2JopuPgSnIdG
FYlP9K7bDmsprmj9clmUqH1l7st33ArjUleY14iamxpinKOJqJFyrfIhnjNz/SA39UklkuRfsvQz
xfLGmf5+FnRGawkzSJcV06tCAVl+N28qFwg/ePE3qyhUl1UXtyu7ZviB4FPsrcq0JrpQuCXJDIgC
JKcQcKLODtNcnw19+VbopOovcynSqv8k3bqhChbWoPUS/IhLpes2BOy40xMKg3wRXDutRloUg4Pr
KE4j1UTWTasFczZ+nWYSA2Oqho4EvDXdJ/BstvQvJ67t4wxR3tgCi7897wgTUNrsFAphgNb1l12j
uAJt3QjKKzSeY26AWY4B2G3wVmAaB0lB3KN4BUi0CxdN01xDmW2UIp/Yvys66/4YJU7I5pAgmMO2
AKhgm7POHVWeMKhIESGPQE5/2HjAh7Xrb6VY0K6jsGTLxfKxXHRL+DXpuOISDranmcY/nboUISP7
6R55A4SkGdScHKbMHXI1JloGKnDmPCywYGVYc+2RyTDcUFew2l82XSKz2kLjTXj+SXpBTdSb0WzV
YbzTOUR9Ur6GXUflPPuTgHrZeMN9QQChXJn8HmSkWeZr4q0LufuwyCR8kJ2CW8LHRzp8E7dXySNU
U/12ny0KtzIflYTSEvCgTB47/m0i2tY2IzMb8mQFblRiUdIIC+NnTJDBOJTsqP5yT90/soPLKyoq
Gs7fFx7rv6/31xg0iLY0IfDVw3Ld/ljkhVOc0GjpMqKCi/ilUHYYb7+BeBMuBY/BT8LPxsSAZ27x
QmGwDtpgjmbM7bNCvfR/z7ttIK1L8HnlgCavqsrOiZ3RTevOXglIQGD1dU6rA79UWXkVknCp6s1g
rpe8XxluH0Ke4xelb5Ya12TYuCuuAkUqpftEoyjwvftEbVnY0fowtQj8SnYhqi7XFWAt5fdAPbKY
0e7WsJkmIhTBTRUf5BNKY4q+q/KmJCT6MRde8zEeKADpDebSEC5CrS3M7oAljrGfWPJivzaG1Wvs
EGjBVLF/UrNxdZuTIwQZt/KUpeCrToxMLrP2auTEIE89SlQbcOEyEGXtNDEphuFr9bQAhFMg+p85
TFc2s8uuAmPfvQwVnMwssFGraSyd581UPu3X0N85HPhqT78RW21kvBGhS+d+W1OlAa4QAajqtFfR
QcLO9bQBZHRQGAyjb3QoWSH1xZOI78eyI1PBLe50dWhUVlsbfm9P/TIM2s4lQjEfEtlFNqmncAUV
PZ0vA9bkus0VcYA/hsrChtWZNT7MOZQ5IfUtNywGvCHh0EXegPa+fWeGEiuOGHdMpkJIUekTFf7+
gT97RemB3Evac8sUfhjjSUzSLyzJaK2ii3l8FrD5cxrrJF8gbVPf2q7mOMT5ZTuAUej995zurfR5
ft9DMxOCzmoCBHUaGiAT45DMGKr2DcOVhYVddbMmGXBX3lL0KR45dSAURwmwvkte/5Wz+nOGHsI0
HY2UXzyXgRx9KWzWKPgVRVrNIXBSRyAmS4uQynWaNdJWrEA7c54wIdyuXCA32Imikag6yBCHcRqQ
b2FnCiXZvM7as1Yc2AiPGG3GEOEkvZsk/azDIsVdfY/x40ousSbTl/teB8gNeRgSOMA3ytwHn4N9
kDfXzySvs/tqgdkrlua9qroiHCRlDffDAr25r04T/o3UCXyH89aIg5WarpR3J3KnEeJnhqSFNmAT
YUhh5XCKJvK/ffYskstQPe6+TyUN48JrciWoq9Da16YYPtooKtIotGbsk0C7yYbiyKLt0cZO+NqC
AkaZt3PfgOna5Nvs1HBDzxeJrAq7jY+xxLsD5QgS/toih4aQ+hB6qbQcmKfWmZUco/bKYVVgXuJa
+RLrEvtEGHLjco56wFQWjxfMP5tSKAIT2a85MpSt+JBM5ze+lHjDaxn4PY+46qydhV0XBEdi3SO+
BtEwb0KqrsAVKVS1YruJsmvm4VjkcdE5WTGOyJFYO+/K+id1bN+E3cjofPtQTazl4UsrYmvaIMm7
kCVA6f8CI3mXh+C+UFWLuae8i+YmVJ1fux34bkWF8fALExiUNDRjXmDDohkdeVKf2sWiQ+sAAv7R
J8QyHFy4a95Qm7BUOIGq4N7ULGSwWn++eeFtCo5o8+M4viugGhfrfOVpCZ23juP5mZ4a6J0xzOic
VopmNfEMouKc/gI2Bb/inbCSHuKNlDvCROEr2Gfy+j2BOeRFgeQYtEmtTA7fY6Frc6H3qdB27Ixu
8gb3vhaQqBcDoJ9ppW3VMIcSGVW/kpLPdx2v5HsgKHpNTj162cK4jKeEFs+37kndyfr54Ife8qQo
XLINFg/dxODKK7btpAH9oudNGXjLR1oZgiygvr+VyXA1btLugG3g+x2cofWn/6sOL0wAFWnLok/O
v8vV7ilhO270wr60fom5Mlx6uTXiFIauSVx2yjZAXZ1YicvzxucC7znLoaTI/q58vFMXXj2kzvdO
tCsik26bPDXOu5gWlC4ExNnFM4JR4qz1zhJ2fagKtT8jhmV1mshPpbo62N+mGG5GBfsQ/pp7ZGRp
XIDo2AUJ57Qf+FRovUUgQVtOb6X3Faafkzkqhvi9HBgl/603anBQE2eoVejSM7RY+vHNR4c0JWiP
3spSjI/UjzXpjYR/N2BoOKB7P3/DIk6kK9Tb7Iya7vHeN5mryHphVfIro3IZmC3Y7X0zpCoA9bzP
Vr6lIWsj1qLiapwwzTViPWwv253hLB7wz9aQLiJLMwjI9vCuW0g9SPZwbh1nH4BURq4MBWLGALgr
In2QovITowkPUxIgAgjFguNTWVIdtY+WLz8XO1wAY8KBqvCi4oZHT3RodgyQ9zmeeJ69fxwXQOkQ
EkdOzcxx9HcYmnsC/ETslONVwvzd0QbZ0XuPk672iK0ppqHRgSUjUaKW1W80AO6LZ9hkokUapo/g
xcnSdJGoOjJ/sJ15KEp+zH+ASB3vMqfx6dhohuH5fEROo5SmAReLcAsVL8gcQcbojR1f0AWURdoh
UmdLvTRkm3Ydcq/u5p3ig7PD8CMAYQXBbXwotTK5rPw1Oq2zHAFs+zaDrnUIXvy3ayK1f1Pbx2pL
JwUOzDBxSLIPFwsvW2qlmEzGKWsuhB4NQK2CP5iaF0u1qhpmoEn0g5Y5K0EOYEL5hAPGN64bxND0
o8MXqiUqofkL+yGNxc9Zym53v5zhZQ0aQRldE3OxgOlCE/63fwCD6JYR2P5CqoQifNYUMnqn3jrk
OT6bYrwV989ljxtXY7EohENvbWJ+t5QiGDq9w0XtE6uFmqZkRDiBNpO65c+Dv37dsvI1AhmlWECr
n12jsihx84VgwEFnfF2s9IQMjPf0kzfA7u1ZgoXrYforShtw0yQGB/MLGe2PakReKUMSlqyxlzYu
Hl7XMDIa/HL2oTt43hWQREugcZ5xOQvQtw0aWIlfSrTNQCIfh7gzfhJb8iLKrq6eAMUGIjjbOsqW
bKR7aL3WcppAinnuypbJkCA4HrwzSXV61w0L0n9eB8yuO/QFH6rWDDIJncR+EMt2fFVcyxp/5rjg
NR5RhnXpuHGlNswqzzYnAP3O6DNXDpzMAuNSPTE4wdCpAcRFx6oxFMo7o1PUbeQ05cNwR/o6+Jjc
loHExYQhdqqzP6Zn6QrUkmHTJ6j1+DCjGA4pXJiPAVvHrNrBoS19SLZb9MYw9oPjs9SUSxxgW1Em
YSOAxQBehtd8+JTDNitQYjJ7V+1aEzesdE0pUMZai+bThNgHrU1fpZpr1/lT6050ZZQJ7PExsEXq
v0AmnPZaZaHTXow/G5Gh8EvYmdFxzMbh+XL8PcDT6aZk4rxyMCMYw0DaBDVHWzIXEOgdQUMZxffa
rq5TXDCm3uNOK2NNllE9UMLcuRbtFvwFj8Hg9CC/Ol59NLMwR3yllWEsUoF+wKVcp4P5uW+0kJuZ
kV5EdSXmXhie3cRs5eZdiH9moVI5qiB7VFVO5krLVjcFpHV0Ed0vDJRiinfTolfbPbQWahMrKna7
UkFJe+FwXW0YtWYi9D9LrivnChrllWDtL1tpKtUEkmr6SNefqfA2OBXMLp16owpGA5xoGEQ9vfPd
q0VKuQg/UQ5BEz0OcstsGanUjpR4ij/NBI7m0HEGXSHxrD+R7n2nRMPqGollG/DGmZHVqZSKihzI
otFWTHAc+kieyT2kiMFhZ0E/CP1YTXoIPsPcWGr3tvxWwv0g0DTHZDXZkDRKBv6WsWTHJPq88fDG
WpCF7A7oKWTxGXKHiUw9YxIP+zQpgVIvdp8LqTfJSKF900a84Fs/T830Dc5FBJpxW3zI79Cj5KyH
EIsp/yyGYXPv8nNmvQVBYw4SOydT0MBqiCW0ECfeLmuGf353v7kJSrDy9aMX5wHGaLnui6/uUXO0
DVvfLOGeTgeuCUGrbJei/9KADHTMHygCcx+x7mjtPObYOzeioh6jZP6Mm/q4i5C17gffAT1/5bVR
2+PB0XnoOoR/J5fOS9JRL3ulswH32LmfvvSd3S/ojZHLR9i1kGDqM1aBe5g9AjbrJIeXM6i+FNin
C+OtQS3z4g1Nd9dIM9jhpjm8t95qbtKykf+5CNAL9SLCLTvSZvScaxA6v2ntRUbfi17XaZpUaE2k
rS5GhqZyYgFKBdamRGDdKCOP7Tc+a+rLsOjY7e5ueRnhw/549E0gYSz60RzPOs1MYaZwstmsXzpA
m15BD4vtAPNRqvewzKZoIk337+9WHl/LTZpRq99UWNzKyE6e9j+C4vrb0hMcSvTTlq3mAtbj5c75
rRFJb8zwE4S5Kpg8cUgbA4klKEjJFzcS76K6Ix6emTDz27RZDKSHjUpp4YrSgaq9y+8RkUcGe7h8
Vjo0FGFb9+d28n0j7Pa822Q62c42PCC9KGNYdNywaSe8IRx0zZJdyTQRxKQnB4PLV/+l+UDH52Ir
yCtQJNGKE/mtOXlubpyqIIsI1APxB7qBkU4hAKrluzR/lI+ZobwtQ83G4g9PNbGnHKRiyUYYDoOt
LOKDUh8VqFlSRnhcyKXtd0Uo4QpnBp/NY58e8aYMI1wnVcY3+OhPksd+LLvpyeqpwjXeuqDTTTzI
hS9IMwDcpTJinzeqgIZ2Gk6dCsKHy/bFv68anb9Xa7Q63VKgSXcB3U2QGGULC9mcZstlY0HZDysH
h+knXUy+SKtauTr8QbGW1upIeobf/+XGewXidb3bpK/fCgvIsi+Fa4SCLWqKAbEBxds0z+kwFCAD
D/gNX1PdW4d07sqRVZpMYCaWenyK88yfZYz54S+fGJRYSsP3GG0qQ8rxqQTnqyGxD6MTxA1OskdJ
KYDrOiBJj6qquKJSo0baGG5WfFb8gpx4/X1P+ZVuA5LWtkOp02vE2UvT3EN9gEYNFTRmEgEtLQPE
9kXp/HhyYLmt1SH6ydtEAcZNziTi2/ZyQtlZ1WDmxAKSQ12G1kevSDKoq9ZcBXMplglqf0eBGB5U
RN+kCjvXObT3aB+rRNoyoHpI/GAlSQ0EJvAAXD1Z6swkQ7V58vSsRq7r4cC8eEE/Fl+NCzhBTSso
mSPLlH/Upzxc0+I9FeTPSafFJ2z5IlByUYTa5qJoZSR0kMkqj6+4foDS4iCAGhw9+I2ddEaNMUsu
x8atapCHq/evfheyd2kxdS4ScIAEjMg9fnRrp3dAj0sk6zQZUS7y9IPTSqvGMXUayoZ4cMczY4A2
dL84cRlbl66ZS55btfXjJx2yExDg4pdB5sF/gFEcbGaK9QNxb9lzzAruzs5Th93wyog6VV6yr0ET
64hLhfD8eu8S+Z0YXS4W4GnhAlpylHatmOfd2/8i19gJgIXH0NRnbUI0FFnRfBwt9hDL9Y+rBapg
IQGmJd3mOkEwhQQvSBgWEViPFjV74ECIoRq3fgYBh68fmQpDyxJl2Be7QIh3vBstFL63jKk0cjkA
rgXea9BQOKm8my6N2QAJuSESbft4OJ4AteRd+j5oBRWwXAV32KVjROx5p2cADT4k6L4sXHjNYIOK
JF8V4WyIAXNx4va9NwxQ9QgPhabIyj0SIZ56FB2DXNdyJXt8sHzoPqxts8DU57F6gKCkJNcTxwuH
rpRx8RISeiaolILsY8FHJLHnnqQscAuM6dHsIbiriVxVR+NDypqPXYfgFo66QifDMcw6gCNDRW5U
yG1GPQ/e07qrHaeB1cTBod5KU4l3DqFUVIifo10Ms9IipY4crFxpBAcNghcJ3OqGw7h1/ZUrJsTv
LTieOJNSTEoJApsJBRPoTx18UW1YvWGYHvSGZzdx5e1IWZhrW4vKerQOv6Yj6DqiBo+Hr5QjrMQc
s2+Kxymk6oY2cpzCkkWdZqOFaQmpw/6OButQXcK6rQOoSiVfZHc5jX1li76eDAJFThgkPXVo/LD9
AHXPCkQGhHMi15AAVJAx2hYIG+kATn5iQRRRi+K/i9MTWAHguM3cFHz5wp40kI9KNqrpwY1zmlsz
cVTY/vJYx/gw49qAjYcsk8o6JeoS8U7+pL+A0vQXdFk46MX3l8L1chdrtZ3pl/zvi6/Kc5tZhzsF
Lk9qJTlcby1K/6v1L36L2KFRL/CQdQYqKVX2+R0SN2KMWReXWTRTnolPUwZfYErqKtKwp1uD4tIb
bFqAEKGpd92A+g7+1rRu0oYuEhR7tWiVr/OKRzbqWJSJXkt3VJ60mJqEK/0zcrYRwbCH74Gth8n6
vMnpJi0pApDtYod+RNEdTxU/P7NoWQCGhf58PfE+myZlW92BIqY1slcyjHuqmFMLaeiGSeiwrdFI
OveRt5rStqbLhopjzYYR7ZY4yo2hwVperQgQkzol4ms+VVIE7QB++0laLAPm3/4ET7F+WcpHn9fh
i3vdbaUXJrtLpfXn73Sqpa2l+TlpGLbwSBytx42lbumgbxxS7QrQqB9hTZ1v2CcwnObY99HN1B8m
z5SxNog5qnC/JgR0EY9B7GPrEk6k3ELbxmoldgn620oLzR/77rgvUubgHuEpyizDVVgDFcuwqhF+
iEpyJs10HRm3zpq2ZvfiR/u/s4iB261+yVJV8GxSzbTZx1JbakVaptMvvsEjj1/Xdm/FRPMpPl3s
wkLjj1x4dnE25GtbR57egscxcUNvSqS+/FvlqeA/WY+qPJrVCPF2j2OWVdDNIlViQ8KMAJJOA3jH
1r672CJ8jzg/xgJgS2t+HIOPQgPQ6/SoIqJ96lLV+ruF9UNzz5ZJmIL94qVpr1xHFFkbuC98gdQ5
C46Bjiklo8OAaA/JoN7KkUTZJ9H75qaCm10gRohnU2rFxY6Lq9bCoAa7eDQpnMCHwiEHAvbHBW1B
eIrKMqS5jyYhnWAZFjL22ErNByZcQMCfqffK1F4YrflIPAptj8r+ePKZIUFurOcDFwRu2mTYLj1Q
PUbNa6ffcx6gwRIY3z5FeLGgxQAAd39NEIGozIHINocj7o4h5Z7iSP0cHQNC/f/bMZrPcEASrR+6
FkuU3qoUSItSoqBrYHr7/h3H2FtFF5bK1qoGWP7ww/D1V13UWFoGJGUjIq4fyTtszeFeBZESG/kE
XH7dZF/IEsPPXrVTM28iTmce99zPPbVfy1Al6dwIEpywg4+d+2ItaQ8M3xRsR1wls6RdRgua1pzL
VBKKwg+QElbyXB3Znr/TwNRoTzK7slOf4LyyFS/yXTXqhTmbiv6pad9795pK0SJFpYfGrcHfDC+J
mBqi8roQKYoNiBpgxe90ORlrs8MMOBLhrNVZunG77K3I8ktOExkUhKJMROZfKcXE1660sg8QOkJ1
08dfjFJ46Zci9gVCU+yrOm2JU53H86ERkoKqAzResgJ37mHZhYLtnC684cHD0NDXq7dHAQBAbWMx
m/xTl9ton6rg/qzWfektEl+DnUmUxPxLNNWhVH2WQM3jJ0NtLA62Z8TYEiGz78Q5Q/jwwtfbfyZI
xOnI7+qFxWaY8qfiIORheE2pj4v0gK7ltoyDo/Q8APU5XgO7+WsZBp1rraJT6+ogxGhvy8Oyt7nz
+HNi864NFN/xBlcQMHdq+qlyYm6BLZOWZbXucydA7o1jUb82CtTDoX7CPylWAyoYj/8u8TA5Z7sl
/0gVnEcjWHMMSOexxKf6AZPfoNWqQOUgVyYaF37ma5sv0yhNfLcPewDZWQJ7K+7OPv9vxKFAnjof
sWI+57LwQfjwOEKZhf9aaC7r0R+D+dmRxeo4lWylNzjFgtoYVZ3G0CnVxdYHpbTA0MWaOEw5n1Uq
QYKhIlZZaozLcGM2OITaSdqcibQGZB4M4Lq2rwOREuigY3uhNn7+44yJEUjdK0ABYSizhE93cz76
8fkaFG17FjMtHrxPWqTUas0d4HkXhIK/b6OpE98LMTNvIYx9OtslTi7F1yKDkma9LPR+PeGw+gLB
LVlFxC07tc5RsMh8xYL7KP3Dgj14CuE6nKsVWHgJqkfS5nyBUjkbdNTuknIG6oFulnHvKV43Yu7Y
jkYp1WxC860FlTlgiXQDhbkKUvfrR4ZbjKNThxu1v9KDs/CBjVQFeasnNt+WO21SDxz0WgnZO9XA
XqNMQlQDnhIRvStspMMd4L6VaTZzrI7kEAEQlvogv04DloZs2gJT6zBrFee+7JOuDFkniToL0wkZ
iya1UmMvhaIc9pwzHIG+PmetfZPYkpkdtOizTlIkXZhheHqCWrHv9HUSWjkUOdK+dX2yCBTP/c57
aFCMzBN/mhvEwvSrBGl3K/9aJVEFOBCyTMagUcajvvnIbIwB9cdtxJafW33yYjlSHwsa3cBky4cN
BJPebsqfZWOKRlCasMQCLHh6NptkdOsY/tEY55cxD6HTC0OWSFEoVkaQyk9hAiGj0JjoJCOc3ctH
PhXqixwEKqTBv/soz+rHgUXLqsYpLOdrdiomFwhDyfb1l5/On4n7oRQxECFVyQwFGSuyLfNTkDW9
kbMLTgZC493Y8rdhwGISAABccb7T7b2ThNLdS5VXsc4yHMh1HeTxZTbg93VvRgp84j6TY1sj42Vx
UXtrvYz+CiW7LcYjWB7aDzkC5BhDiIcVluefipKncyjfORPZA5GwgPbdf0yupc25lVbXHz5i+xGN
sOo79XfRbL1KJrD61P2Rd/M3mtnxIYqQxTek6DRyUT2fJVZ/AWc06MiND0TnHvl+c3+W+naGKpiU
y8LcZ1WvGvC60cJ0gD15yP5adM7mpOB4nqrjo8BqXzLuNRaGq+WS/x39MYt23oaebOltZUvr8kCv
Ma6rXNjgOPDGiEsdx1zJd8Saa5GQq+mfJUry//Ew2KW9JZtOjlfmzgMJeMmlK5g+eAFbt34hoxo9
v+Y8DOebFrvPvTFFIJV9f/EYwnen97jq7zjMCF4SPTjS7nsrB3mM2RwtQMx7VjJAk+6DVBXKp0mI
mI54wu2m2uIH2tcidkioJCTEDoNCGn4op34TyUt1Mhk/J1L80Pmn6AE5jiGr7sdXaBkb8L9wJTFe
KE8Nf3e+viKWduVx2qKNtpyeUdpUidccBUnh7TIswBzEUv+GLrMz/PHmpSefYp2nZgLavGAm8Yn8
82Qy4s6x0yOVy2qFt43P2BODBRv5SXpro2EuQM0+X3f1C/9liGdBKLt0H6WheptnM2SBO3Aa95nR
y0cuntWGhpEpyNhuusmN7g4o/xCOzOWHei2DH0DdjbYXFUIuMHPEjByvputKmBHxr51j8b2Y9M0Q
rvjGol2Edj+ReDGwFBCFSRq/vNsDzpP7H+/cDyrxaTlfEznb0Vi2pHkv8qQBULPBtmrTOYCo0JVG
spbYT3/AbkPYsyFCGYwKTCNzfCqyhnSlxJCOC/q0syGk/R9+HCjx0v62/Asl53XIgxiYGLU29v3z
wO8MVtdUH73BHETBvMwl43FYVVhPge8lYGBmkI9vh+I1TJq5xabp9JwmdvOUJz5QsWEACATBWXyw
ddohpp7EWCT9E4wGyJ4vIo2Qb7CCOyO5YCzVPo8yNtbFZLnNcQTdKof7lHPbXqXtkrUrTMiL6foq
djiRe8ILM+HfXe7mkO5UIrGzVYY+vNe9NvBi1vXNmvK8VJ7X/H2RCtryTgmrg73AWHACuB4iBNX4
gpcBUDtHp2NMVaTb0CvEC9FeUioye185ueJ+4R4Xc7DGMN1OLVySm53BiFwGtMVpHi0N3T066omq
oqzjw/31NG1PVrBoQ3EbSIZc4o98ygHYOh140zF8yLc1ZIsXSqr3pZcG1NIknjDArRO2TS1I6oko
Js7E9UFRhzOXmIXoscHpeI10jlnVY/pHskwe1Ot61r/u9/A6TQ94L2bUNgXkHZpJgxX1d0U3X3BZ
NRbckEW4TyIXK3BC2R4ZgTXHqVcrSWGXwXClxJuvrW0o9Rfr5mrneNi2HNx/GS6SsS8PEoUZkDi7
Kg05Urz62q2oNPZqyFuK+GcevrvmvSbVOQ7wAR62/Ywar8zGW38F5n+np59NurJlXlQ5eOY6KAlQ
85GYqfcXYBFDbtMqdqYPprVYsLJs6s7EMNCaL/IXpdiff4iRXbE7GlafMLpLjhr8f65lQSmduX+K
maFS43V9T9FhbdKhFymGNdYOrUkFjN7CKvnecrwvD9xwXx55+uM23KdjSUpaB7fMAotp4qwro9OU
Mx0e+rXASaXcxqICekQaItyWr0NzJRA5NZZLLEa32VqPP/+c6Amt9v/j1uM1mp4NXLNB1FvYZAIV
7I0vJJM0Dvb74Agy/bRnIbox1K4nouYYvYftinKLUEYP3CDdXFhwL5RvymgI2GoSGg+VABrq+UD2
f08DbhQQb17dQbQa565lIIGB9JCyMvREbUFJCrxr3aEthnLNF4wEI01+cYj19VtN17NsRiFP+cKI
fgBlfLsR7oxP4wyw1FGoH9UUOCIt4WmVTb6NdW/cix7UPnlP8OmjdFCXOkOXlSSY/eOEbCk6bpi1
Iu/0gVXzak2fDeHub5E8+0P8xT7f0Lt1S1F2tp+nk9kDLQ+X9yh1j0jr9lRMc3WXxUZEz9da0Nfq
Xift878N5stSc59QJ8LCaOmg6dwWp4E93sKF0GFqY81MXB7ZxYyiemCcE0UDOpgSOCgEhbyai5Jd
PCrTvP14c00XNoHWyT+6UdNcPvWIxlzhfm2Qo5cIr1gie70Zbqf1sj6ENacURLKnwIuf2O1uuoRv
FdxLRBiUhpgweb/0GP9W0EFz9Hed3IvJ3pMzZzBSVV5E6M8bxmL/A3d+ecqXJQP+lt9T8YhSsrCm
ffLV2M0vg8aZgxDh7NzXG1b+u2kHx7A0wP+cdAcGxWEUsLcz359mp6GBrOOVVmQd29HqM8qaCIdG
XkUEs6S8gV8nCaGd8RAxpEygFxvXY91VyFWD47vDF0qYZ8RV1N/kycdBZN0o4YO8dJbFHGB4jlus
sN4VtWAz8quzjUuVtqCsKnbmceKeAho/u1Ejb6pgjJEXUfjd37FWLvYRA0aYM9W8AVu9ZsCP7Phl
hYUpRkLsy8BYnubdjx497zb3YNcePcU2zQ0irdosu65hJa4JR/8SKKNXwURz2aRani+2CAgGy1Xm
hpq4+BiMrVM+eXpD0oiSbBhSsESr1NGTzt3zeWqAmvkQcddSaKvTFizYU3Wv1cyVClBFAd+xhL3t
TqyET7pbhTPPmhte7SSFtLZyNAOeBiZxSRu4c/EPS1mIgDm7bwIoeX+GMr6kv4FJTwP4z8wRfd8a
RO0JQpjFlhzrdbIqLyMEJkL04aTlIbUHACpFQEHuX9XqLOtSMvcW7jsEnJxtTbc8VrIifR/4AbAZ
/M/0AB5Fz2jG4WvwRAsBOmV8jTKh9tgstRS7CxaL1oXocKAIgMuZHanINHHLnDZ17wn3AgvGxtey
Ow1ieB9sZo0qu8ic3V2x7BKlsdvPnRLPeyoNb6xebbHJPRIv4iv4/HmUaxvd9euB5NT0uiLi8ZM9
SgPMS4nC0kxzheZrdmFH96a+qSNb0WjJS8Geu281OBQ348OdV4iEuUqsqBKPiORC6uGoy8WyB69W
EN0A5ODDCKWBHQw+S5kVwyZNJJYwrgL/VVkRhqhIT3RMiK0EG4vP1e8YII4SEsq6q5I1SYT399nA
Gde1O/Gj5gfoEaQoGRkf9GYNweV4R+N+OzQmQuP2TgppkSOXOQvT/YAvxBibFA56J8k6C6Xpin1M
/XejbAPxrBexP8GGb/NiC8Ekd5EwZ8SBZBcjYYsMjKE6JhgjuSGa0CKqpPLNrml+mZVCTlowWxd8
plQfD9iiuj4hZrLd+3H382MTZrgJVm0DAfPi/+4N0ftKPOlPNcRwo7afJ76D+qRLhPkhJWFCk0qa
q+9kImhcQSdUcHzO8JLaad5E/hhlP7bfoto/0N4J9mQZLBhB9BdJdl7f9LrgqJ+T+6Uu0VJuY9Jt
/JA29lJgdx4QDSPIgjulSnQAHs28vtShMogg3Nhv8vcTRQgT5kVNIsx1bpi0TU8VjCEBn86+semC
Ey2uadN6ATKOtFbzuqfQOgdH+DbBfUhUQLDEY+co+ScV1YgzLPpiVuN0jCBNihxdsU2GIoXZkNC/
pJqLXfTPt+3lVMtuxrncybschTZFpuDU82RcRs/fsn0ROte47XLaA/bvAIcI0t65qIfuYaKfKE3z
3Zf277M8rMHOrZkHDIJR+hIOWohpWVrMM6lSyzQSdsnEffYp07MTIYnUCGcP1AlbVf5TNWaba6et
d3EyiJxyn3stAN7+9Hz6mfw/R8oBVbmwNJbe7hoFpUfF2IJrA1Iogq/EnYOklZxUMC8ZDmQjvTuw
b8+2Acip4eDWgmRyy70EZygb94KP8xCODR85+N+ZCQ+nS3ZmPDmZdRfuFKO4KLKbAgGGgC2Ypl2e
+PDFib6pcHM1j7Hilr0kNTskqmBthlPZCR3sa/cG6Mvos6qUEw2OxFjWYA99w7y4jI4XId7HJQPZ
Ve7Z+x5amnGSFsrp1NUcSzw5BkNfvNfSlhGH47ucfvCfBWErIEB/qm/WNTIp05xGDKsbmIeP64mH
Z2+u5TyLjHi5ko3UXLHKvini0oRd81RyLmKr9qf/ogu3jnq66SZNouGlQGjKmA61w3+onaSvZP+B
2zrW9FEDgz9cL95NYCAcXtWrzntBhwpu6tx0pOLkQb97ltjr2jMSDKIqe/iFQ0IWGJL8/V0cqscV
y2nfezcwcuQrjmOrVfDSV30eu8uq0iArcFw1wsmjKgwrpOK0j1sN4Cl6FxV66dB6mEi2qzvDRf2V
RhKnytn00NuAjiCuPAbGVPTmEmgyZZtaxivZfRST6TSByyOYOYEOa69TOjs/nSYr71LimyO6ZpSi
8/tiBmmNbGRAmY08eY5ayIq7tUKoIhTKM1uIlm34sFeXcYNMHGnu6uHZ4DUKo/VAq3sIpR0P66x8
zaaRQGa9QHq8C01wfQnptgGFu1w3QouNUFcoWGZDDcFOLLuFXn/Pmew2PTWAqGY2qNNqtPVm2HiW
FpEWHbcTbI8EUg/QxnDhuX3dDxiVYbWvlnnC95KMSKvT1ZDmXq8VBJcmxgK7Usir0+lpaBue6dh2
1mdz5d3y5+PEpJa3TQdI3cnCo0EInlUkAyf8EmjuzKBDrlS2XhdS+7aIfQM8lauBL+evFbV9uZb1
AKpFxhNoyrvcCwKUcN5+s4WmlYViLf2dkqSoM5COx/mLNR1+lrOe5fSFmNdrijOhfvNNyYStexxY
swPusSCVyVUKjm9tFNb+B4iqg8ykvNR11k5vdUN2Qq8ts4zT+iJgUZCU2FDP/ePl4Yu7uYBJOa26
KxaBXO+RB8eVqBzGSBFqb9XSjRjdqPZPOXw+VghlyxhQuRbMt+ctrmgGH+j/XHQprzpiNJiih9t1
s6eoJ7t6/Y4yJbJWWl2imW6vczU88X8ipPLfu82faTxKzapayh4nWgjMMDi8P6htqpgmTopmo9LW
6NSGuUL2PVMXHv7UYIAZPjUhZodz1r6XMyscG4Jot46qJz6jJcmtgR+M3o90W9GIjqJWIbqegLFQ
T49l10cJc0+c0x5Qnx5N9CWgt+zN0EQX715zgCPVfg/rNw1TvTER+13WqqI/amIyOdw6ct5WCJap
XeRCuXDF8xaYtzRKQVxFiAFizJEyptjBMJIdkHRy/GFFtGvUz8JUUwXUpKXhONlJQ0dFH2CY9agn
KRjGvydC06V5zdaJ1KCHtDMpgNlRtusXySsV93rB5d8cpGae/8xYmFB9vqMktwrudacCa5Xklxrf
T+Ko52ePhfR9paSFU6PW259Pm9kuSqZE9K+99+6I6VzSPl5JZ1lcx6g0VBiDueZA9h+IByl6dvlO
rHsyNug6SDKdeujemgIfpR9/UcZzxJmNta0NzTEPanV4UZwiMcPH+ER7ujuARkQuuLqHXuVpYTvd
gLpQzoBNUTkxNNu1dOM6qvK32QI9vb8IKjz0mU93kF+D0pzmLfomhYG/33W7KJWFMNPkVfTlkziy
3SeT4wJ/rZoz7dn3hsIPHlvrSIrvoMsKXyFL73zOF7MSjYcPaBBi36jibB51sqOsgyBTNE5i6tDL
jfEigf4F24wuHgeWxQGbRlozY6y/YSENxe80PiIuROVDWHPMLwpt6W3tvLvCthUEl/VKxKJgITcu
YBvPu4pHMBXq0J/xd/JKXTCCPUb1edrhQrctLnDe34rLIThKd8PNyT7dXUVvou5j2qMwy3WZpqGu
6oUa8RBLlKIkr7yud4lBphXGYSFHr8vF841TJIhhHxFVPjA48gXJiY66eXD6cJDLua/GakjlQJ2S
r08AWzboucy1I+CQaEYcuxxFvWkPGRUtf/Iqw7y11maeNIDgxjqIhvjQmjIZt/ZtreYZGEHRGSe4
xHsigkxVbqExrFkjmqj+B7/LqwdvvF2HvORTf5yufIrCPmXwliWu5uTMNqLKU1utbQlYQikMwC9G
/KRMTBAl3oUm9yuJOfSWI55DoKOI6fp7FQKeZWLmMtWJDWhDhgrNax7q6W1JqHwhkCj1+vGtm93e
BVtF/IPFiBNinaonU3hrT2l2IJvK+d171Sm6WB1LrLVHTcx5ftZwC31IY6RBDL74OtamtZx5Xha/
Rsky8eS6Xpg/UVLSHp30IwjPipoaB76W5LxzVaMb0ZiDALWTeIG3TysflEnCeHC7zmLCbGiYJ1nt
Hko55JWyalkLOnRGyf9WdLJE+5LC99aNxeBlnkSXohNeoAUC6RGZHYl4L+hna+MnZRZ/lFFrAeFZ
vUuVpKG76WsRxKv4f++JHCteNbl2gBWUtmgQLo0Qhafk8Xc7johBAPWdeP56UftoKOI0gVXpQogq
qLEuVefuvJpJ5/Yod0kCWZNdvoFe8yx79KCQMxBVmT5LN2H4ppI8OFGpeUV2O60hNYrkpat3H3O9
rRdqu70eXBaUgd8C/n21P6YYLGXMq6QxEvE/67fWp3Q9n/Rnwkg8B7D07UwvoJv1iKwUbOWPd3u7
wwY8NBQF/chQcdsS0Fe2eDbbqdyQFZbWvkiD+eSt8Ekag89vUge3XJbfq3VPe5Oz3MVsqSpEjH/p
mWKqCeb4Onb7404mqj2XJrnmsdNrtDulF6onfH849C6tQDylwvgmi/87FR7dWFgj58Ky0CzbsWa0
2hZq2ppdjWiJy9HJF5yt62GwROjj1T+cbJHd3l+ox/DwnlLDbggNm7UPlXUWimCdZ2TGTh4IETGo
vlZNxWPIWmiYf3zlvhOWFodNXHAnQUlMG6dexsObTq0qTOzg8kgFMwqCJJlXE8CteUKotAWXKyxg
69v7ZhSclwtlNnX1gtJT6++uS8oIoavH38mOJ0H06EkpEvs06BnKKisMb+6xNVMuQSBv95xiQg1a
zHQvNhYfiMgW5U6JtDbH2wovqh+JPuAUaYsVdj/EBcNJ7AznB6OAoSVgDCbkhHigR8hh/aWdfUef
qAd3wl6WmZD2q4N/FJf4Hqa1GTuUoi47nS7U3f2vSJ3xEeS9jZjl3W1mElp3x/hGvfLCivt5tW/Z
4GNiKE6PL4K+duKUUBda8MptEQnVTct8OTMLLTdZ/G3DvGclS584mwquHtWm9MtT23GOcHyR4UOs
OCgZMrySBLKJ6vu54r7gFTMdT9oqzQtYli1HSVOES8D7fIb1XLDm32pNM5E/prZ1jrZVFjEgSbJJ
9zMt740c+dBpnS1b4l4uKwxalfu0qiGdAmjx0A/vi3LREVDhIuQI2O0izIa/mnXIfZwBGQbqFGHq
bB5xqda4C1gG7x/1pqSrC4a4fXoWVSL3Jx+GMYKrM8jnqNw81qoIaOa+u1mfB1iXI/x2dz3s1zYQ
gfy2PUQG7h4vfooR9rcG6cujnAlkKaZ1OhjCG3LYQtLpqeW5fwusqFHE+bnOfEd1B10NjfPPx6UX
cqHbKf41Sart9xRteVpwXcVvxsRmMTiixy4zLoXIXzsxmzxiYpmujAV+H273F6yCWDRwelgPIPs1
M83WWx8coleTcPcnPgDsiYICE4DeRc9yuk0/dc3Xsu25y5pEK6OHTS1Qn4DHI3vaaBG+DFTH5Zs4
HMpIb7iwtQC7HrlRdmeIum/qq8W+Punua8nhCAQ+Deq28ny7+slGBL7wXgbqhdDYgfNAE0gSPQ1Z
WO5WUryMYDdinPOUOuKOlJyr8dSxay77BpXCkX0Hj9mDeQoNC2X5DCf8wtfsEW79w4qkzo91Q3Lw
f9lrG3r559xW/9xfCDwCGpZ0CTX20oJ5wqB8fRGIkzFi7ibsKRcUcJ2sdCjK1FcSEqa8rO4wvIcH
HpKQZuTvZkfFNuhaHJvO+KdSNzPqpSERCZjpAbayVfC5QFRGQROVTCmLX1TSrQd2H9irc+cKcsuW
pgntuS8aitNr0ostBWUWEwLIyEFAFFR4JuAKp564w0S76gCCdjG+8Vt+vrcoqGD6HSN66FaArtMj
+OnmYzljXKigitFBT09XJoBSvfWhopE3XbRyTg5JTKWiIkA/YSAJjtCcqMKVLFpQnyGEZly5cXJp
UnZkZDqJAMk7syWtvPOZ+ycZS0fCRGvq6dPY8nGgMLYZugXECetsi7YjmQGf8YcZUpFiT23rNBR2
g5DwhZ2C5AaRMNhfeF2sTygFTE9xs5yjowtbic70aCtz5uZHPIwUksxK7H72MU1/xXt9QJRbgvYB
ADRnOp5JLRcZLb4AuTb/9Cm6oDApYU0LC5ReeWcizv7GbZZD7KJaRzG7s+S8s1y5mOmPl2WYn9Dv
R3XWX88RWnuaEmbfvolts5iB+YVwRhgk4Yqfd1GarRmsL0fo6ksTKpcxg+fkMocKwXqeNdEXsSdZ
HpwzDDvQBWa+bGBjT0jnmq94CGcqs0cxnK/Va2DOP1p5arHvai1D1IZuCzKvPE0LYikolxbWxu1u
AULAeAkAU1nlouuJcKvoFgvjKKtX3yYoP/aZrcsCfEqN0XSvi38dRnG9ZiPNLHx46f+x0ji4n95u
s+3+QlvqZoemTV5Qv52fjkUcPFeL8MEekggkqEOkKq6qFCDbeDVl/WBCqZgTam178JjYXeZsm7Pu
tOfmLIAlB3lkPdzjMc1iKj4vnYQyOVqyTkVFsReNhd/rgvgnFeOcQ/UChDTiV8SEXMPbiZfxvwyg
7zCkOHIe9cBwBqBt5g/HQuzBWSMpnHh2thH9CdiIuxh255QyielODedFAzrxYwWOksGKQ1tHMcxE
LvHz2JJ0534BC8kPKMpG9tY+PCtMjRyLUdXbxdRTrXOnq3DIhipE7vHZTITgUpopB/HjSFxzQT2r
VszefQJua9M76jOsjTroosDJ8H2d5Wtj4txbRwpn+ZohsYmCU5vCSTOGfX6oEVmV3+BbHtFiJVkV
jScWrzZTMDv7Kz4SRSFUArmr3E41yNCtkzB3KkhbDdZy7MCxTuWCLDVqYqlgf2n1GEy1uisb3tq2
4fwxVSUQ1W61/gNRt0ECET5fqx49Di8PV076o3NBSdb9h1U6Srgf2Vi5QVXqfwreO+qLYNcKmCgW
KaUGdiZa/y3N/lzS99SeKz7hr7H2AkL5i0Dmf+g417cP1pcR0LeIYCQkQgvCqItTWTd91+SKdK8D
ehk0XtJE4Ol1nsOIKD/SdOOwwGkw3QX39DJlEt/ZjIgz3g1ZBYTFOpbQbOfmoEyt3cJzERj3J+K6
gmpiQ4Bt7XjaEbagFQeLSzcfxMzJovr4tAS9iGtn8luiJohBk1kDPaX6uPJxYFF3Hn3Dj8EWEXne
4keCnWujpRJ+g6mDmOJyTgmUyHx/qs0x7wkaF8qf5eKZKU3czA4MpeBlkBrORjjmLxer/l8P8CzJ
CZk776AzFjWd4uTu/83Ir26KfE+/EdUpgsL08gtUEplNxwu/mf4ZN3T9EtIOa7L9RnvRJ6az1WqL
OyON7Yx5OP7KyD6wpue1LwwFg/zUoBiWnlL/JXiYnuRX7utYDe7n7Er3gZW2gbHodpaYHDdXDKoU
FVQbGxIE5H3f0hDf5lmTDkV1RLu0ePS7snjex+BorYM8mZfrj6MBaoK8Tynj6z/Y7tk5IIz4IHC9
0w3zsjidJ+TA9kfdtOnQK/SnUSyiQUPCrM01JrfOWuJFJ61Qk9tht0cQc6YktyaTZSQnBxCPRf2e
9aUEQh0TOwq9GLa8iXBpfNCleaAs3gdRX6aBWYVWAyTrGSd5POkFwPAI5E8GfsiCgnx5lcPV9O3m
wZ8RfeESWFeCoBaPSSoc6rJ6jfZgKeeorPczLf+l31jYuXZIk+mo1G4a1xfX8Nr36G21qrt7aGYQ
+x9w89WCCHspoPhH3Tq/t847NhfZ6UPmbIx9b3RVhtTMzohf0cP4CGBAFTC14VSOzCKbgQfkI8j5
6Bzfkol5JmLunlt54T0mxTiLxH5rffrKRVXM1+wdt9+wQ7yePD3pc/xH4yFv8bWfI6Kc7JJnEHBt
GdPJPlcahW6K7qyvvHX6RkRv+imMjY/+6c6CIGx4OxKxv6b3for/1lBBs5CmTMaHsV1rTkW2Qw+W
QAq/7/iLHUxg0vGAmeHPyI15T2KAGK0apau01BnW5l3uMkMQB0oADTNyIKFt6pNFTFosiiVHC7zP
eG8NbufwZ2C15t8wUmOrkjQVgrpGX/uiFjRQxFqv3vq3DcsR1qXjj+G8lO6SKjSkZs8gxBhSLTSj
pSBuJgJUx/nRrOcDpiy/p9wBncW4OhffBD+/Tzps0vUsO4t5T8hrWRc6xc+dX7rH6nX/ixTmfVdB
M00l0nkQT9xe3HoNguVb1cNHR+Z6mMw4V3HlxlmL8iJYFNE6bXWqI29XTDER+kXpcxctfbUhAmoG
J3G+VOSbPtOt+Ohoch6Dy68C9htDQ+xyYtjddwZf7CQsWbM8wvHyOHc1TdBdeiWY1jNA2xMZAvIw
FYPGvHQZYxDOD/b0/DV9FVRpLYAhA0qDm/LRsLvFXOC7eFBGDYj6AEReQ1NIb+x0HLe+AaNd+t1I
jQQJuLJYLbeOZPQpdxRggY1RVHNnvV13MQWu5XVE0JHlXC2W1ILIN0FgngFsFn2aZ0x2DZ1897Sp
Q3li7lTnBEOVtMR4sXJKzmbI3f0xn4Ujy88cVCrGqgj+DQi2gl0tGnip+hU4YZ7Eq6MO2BpAnrVF
HECxQP6Oq43FDMNoQ8fBXvDGALjDYcudEpQyDr17lnm3IC5B2HFiGNXtiZ45eiqFbExA6+4qHpsD
uiOX5rI6uSo+bEdXb+RGIMvi5in1CJw7i7VWm4Rj8dHn6AcxlrVQiFVV1TdLcPQ/l05DYmqnjI93
UL0tzwnAZNCnVoRX7nz8seFav+c4vQiZQr2xSFHpU4xrczddgQBsbwDPJs7U67PnN+l3HgYKCr04
DBA4CPDq4sPvugtl/vCfB2kMeZQ9bg6vxlqcoQPkFTu6xnSGW/x1YuWPAwgCVrBANkmUVkV9nrKA
cvxfMGKJJPvDkY4pxo5q3I+A/pVEWTsy1GJ/+MnWh5Daii3F57MWNQRtWl5hW3nS6Zz9imsNhhTI
pglB99p78o8xnzIMTlR+TDJhftXdOs+nbjZQMBuGn/ODkYLn2j5K9HOkPEe3DEaInDZasXaV0l1V
MGoO1JABEBH3lVQm9YerXjqPk3i9LRY7iAzPnay89cyhf8c9rvqiqGIC2J2h5pLMjapejvfEg5/x
ifeoOC+tjpW048d5xXkGx16uQRJhi3jdWtEaF1/L3mMz57ftzy2NBolTqXRBLf7rK8sB3DIW4kHW
Fs517pRpw33I63Iy677JV1KZNrl8f9ilsH8bE+t56Ez+NukMqzVN9dSPg1cyt3Li+QrRj1yPIQJy
PhgT5tepcpP8r95CKfOQgv1GzC0kjOLfzm+mlAeKRC4gGs4BD7yNlBUh+Ss5/nfh5l5X1dbTKgSQ
SRY9CsMBdbqNDrevigpxwo1lg49RZ0/9W4kXFkr9tP3xWn0mFuRVZGbXgklguHkDqMjb9ga/qeEl
Go/rEbuyEkf2C9jmt4nu6vLfcwu5psJoJb93hqyGRkDqn2FlJgdt97Bi/NGMRspcnOF35kSF+ssw
jNAdzC6cI5b3+WIB6dLIme42SOAj2hvvcldbKYqORctM43NOSfymCF1jfNQsX6NZCPSenZ0XtRzF
amfyeY8GQXDYIOpTI8LiWJjQKY3BB+R0kTA7MRNvILR2AFcpYwMxiHQtzacINzGHEf6R6Zsy/ibc
tylhjnmClY5/Ysc5Dv3nvX4d2fG4bSdVSTMORWfpJL3dbeMIWy5EWtWC9nTGffhVGiReFHGfxR/C
wt0JvvTD6FLmFF/NvZQ42J206X76SPKcfvQMhbTk/2B7KNTManOECf0uzwDh273Ibi+Jr4gVe3WI
SSnu5f5o4yRE3NDPpP0lmZUsvwk9i10P4mn35FhMJcvsCD3k/GkMPn1Woutw4VY17vU25WUh7TtX
IIOnujYHUYYkAHIr93g9rLn5l54SPYmdPyZ2xe8NIzmSnBNyuLbqXfy6ziY0F5Zl4nvq+EVSKM4N
BL/slV1yB9fBsVKM+YbLOQQb3tblDnXoXKS7zsG5h/Rv/3Hs49dVeqW71lWOSVZNuei/M4xQqe6w
ZuTaEjOrHJnjh72rYNAYMxND9sVi+n0OOv6NFK/9FDmN69d/jiQ9MM4qE98up6dbkfBgJynz4dJH
i0tHOjljUIjH8AZXqXrkLFyJ99vWWanqdtWkwO96GcUTum/U1o9O8a27uekj9FX3j0z5GI6E8vRL
+o9/u+F2c/3rul/ZQvDb3KQsVw4ITt6m4TGmsHzyc7vPUsCJknSTToYo/U5P5Uo/VJZNkKToa1RW
+rhkNrS8jAe/j3VGsA87wAw1LahBLxIjVanwmDGm6qCdhyqCagVHD9FsTWEYVCq4377T7MK+dNpr
yZHO74vtqPRxAcdIsaSrFaz+nvKrjkz6Nak8UD7MZBIRRSpFbnp4HT4DjDBB4Iy5FRCIW5OLh09C
nzXaZfAeFaGw2ITgiHgVJt3+vLVlK57g6SBfCZjJfZBv2bU2LI7KkZZ9oZxDoBafU9OvfrVU4EPm
Tu7mJAxcaHctnqaGqmoFC/Ds+c7Dly54pKoeSVOzu2kpLA6yFFLxV/xNejwWZX48xJfJCjuxrUz1
Ps84PJYPKmpY8sXLNvRSZ//mNlTitbJvszP7gsN6jqcD8xEcbVnXzbY5w7JVgy6pGUsyPsm9ue7/
xCuLWal9ppq2au2ifMBlpe+jaomhF53pQxtplMwfliSwqNSIvaNdv8gG2foyVsdb0o0RPYbd+hTP
9KHVhhz/kNEpl17wrLuFBCExzw1N442461AF+CDIo0gsGTOOQXW1Bka81wynnP6ojf7f9Dbwtm1w
UAZya1B56TXgE6z+yP9OtAbqrqWCUrsOr6Rfuez3ROtxbjMATuUCGhaLmpfmKLG1Ii/S0EoQskYK
bOCDSDyuv8S7BlcthMpr3Ms+hduz3YF/OYXvYyyPqtT/co1iGNqR5suE3Wg9eYGYwjYZ4AYZZjri
74ay2Qzrl3yTo6zaesWZye7OxZrv4moc7bjAzGOfToBJcV5RWcQKhoLSn2hKVcdyLqT9Cwdn398R
D2uJootmgEWMHgZDfa7ckOOyT4kDfDi5Bj/VTY/tvycBvpD82XjF3KhK2zjussRnVy9RWd8qI5D2
v/Z/VpHdWznrFP+6IrOK3RvxOBOh+raKyU4IZuBdoW3hP7xk3XT6i/FwkKQqT4pIdPvsdSLkOFki
AbtRs/3ycGq4TpW5xjafj1lySQKbmtr2gR0gRsOkqLK8n0m4mtyx1QW0luc0P2AbF1e6gfD9RALy
j13eJq86y7r1cNJYf9ASgCHyYhdw7PhI7oNyPgvMkOruydk7l4fGn5ExnaqL1Dd2w5Aom4UV7q3k
KvJ+OPjuisAxOLZWE6XcJyu97pwqwwV2yIH9Zdu1DZPBOH5jqcFtbgSTeHqBzThuhu8j0iR/XQc4
QnN41WUwltAmalqSlOAm9lpkod0Fh45iAexdrYQ9IXzkSuS4jWlcnxlHHnFnDCU7++CA/NEW7Ble
XOdGdrcq5sHw7hhVJEhUXvvaQvL23A8A/wRoMZ6rvOJyOohIQZacUJvSxk1aJODkt9tb/nA1sJuf
9QoBMJfZLYunC4+Q2EUXjmG7xYVj8k0jraBCgTPbJAskmEM9ZfqEM12Ly34o84qHgXCwynkmVI9I
iMKXXlthQosm1A5GZmWMbToviIJBB+nAdEOai1ntvhklBuHpv8SwvvuDQfwhHKI3zohoIpO0XZv5
AG0+IhnRq9fpUeJF9AyXmqvHTWdWoHPEpXnVXfay0hbWlB/rVpiP+Jl3HgP7ZDR0Zu1ZPBpenIrP
EG6eGH5UDgdHfaeyd7WiGO67hbaZamgoGUV6N9BflevWpwJ8AYylgCbKZIYqRouRUXQEok6Gezil
uknY6S7i7pcZFOZPKPPsuFqRz82jajVL9PlMy72Rpj/TskZ1riTIrTq8bnutwzqquqEXU0dEixGU
EiimfAoK7vJtdUEdmb3V8mISiDvm3QJYILqOkkPnw98vrqPXjU0RFXVRmSY0rkmd/o+VFb6O0kD9
eS0PGzvPwcUyRW1HJl6dTh4Y0pX91iTTIKRvAQxxQ8xaRqsnuwi7rl2IbEq2gDI3/3TUemztgDZB
MYh3Vn/CQCpxVJPTJfUlLxt5y0LuYxA8A3W65ra4jbVy4b+8bqWAwKm0Ff0g8AFbjWfWXXMZr53H
j+Z+qaFvi+doY5pX4wOhfTi5j/WdREzXQj5Seqc0NNMfAAJ8JxmPE0yotR1NpD3unwX2a4hAD6J8
gxAeGvJcPHUpL0IdREvrTsjmj6jgt9/Za1NGP43cpp1usHd+hBZz00ie6iI3+pZ4QvjQYRq9uTXH
nykcE4YWXy2J5/md1YXcloOOXKaptYdrVQkg9p2a3UjNFT2fb6n+dBXTbPzjEniLVVM77i8TCpdz
Z+Aw0emhq65n5pk0DM1WmL+TT96xdA4lV0Khrug/ycQe7l2X0jWOhJnHTDTdFSvu+ak1+iA6Qmq4
TjT6yL6DNF6GTWP2YjxDqJv/pp94YAruHV/smtDYKLajtxcz56kw99lxGxA8YUPnkAw1YA8lLZ/j
3bED/Gmhr1Xfi8fYchg4SYV/eZ75IUIIi2ma3mBPutTT40Gj+k3dPrCoym/uTUI544X4mYHtH8+9
4Ok6fX9Nzvf24Vo9VytKPYvtgq2Ic3qvge6i8L3zBNRbohA0mTCW5qr8rMrcx9+o+gEv7VMUrjz/
/x4M9BMEmdS5Yp9VlJtKr8m4kntlfTiuW6f79EAUCREwkZB+KPiWKozrY2+OcPdThUpBacrzrC1e
oPhmsaRqUwYVTaKvMzhTa/nlshNKHYLsE68CqKj/pwi8z2oHDTAVRb+OiCfQuJGgbu096doKeXEJ
c9lTjB9dPi8BP0zKTsZKOi5I8j/pPnjvhfc0P7xGC+85h3c419jc2q3uT6cmjGRibprCKXo9EJFx
fmomil+C0r+OJO8LnqLG4aSZ3uUB45eOOM2mIUnaE4j7v/HO5rqZ4os5ikUBNJDP8ZCqlbbgcdP6
3akiGvVVx/eZiuirRgfxxZ3LAVkb9ui8YuReXj2ViVbL8Gpsr1s+bO6m59eleN59Wmw3CUTh5dOh
9mfXixdP6PXSyIJPXFBCMx3n0GyErQk9TM/PlZpjjd3kj+NEaKWV/Zd7YzSznKHeprpU3RLf1HpD
MCDr9/4JyKFmXXqmcuqNDiY0nAbfsaswpOaLDfUnf1BuzKo0arIK00HD/PDkOeoJ6Gikug4gG+IC
a5rjuA42VjH5t2j49fKgnYMXwN0/uYbzJzXK6ZZNPysSi7dzBnjsBQePGb+KeRtdJhnGiZFKXcih
Rwwy4S+yNKi0JgGqkrioFygVS8q2VcUhVXsBaVSZ1AJrikYurTYZA1a6Jqt6ANrl8sSTjkW9U3gp
HqdxkducP1q+r3Jx2rdNG2L0AeC6YQJ77mfwdxIOzwOvg3KMzmnJMWXKuEQQWVHetPQhDSy+ESt1
sQE6VKDSbfF8LgSsnB18jqcBT/m+1BxmtDIzTWtrK2fiW9zQCNGVaU9EjZwbWybBHKiaXn/Crp3e
2fnpGliiMVaYCiMz7zLb3g5rzbOd0BsODddCkb4xFtMJTwZa24D4blUfLJLLAwlwyDkFVh/2LNwH
pWs9cmIx8C/hhGDk0g1j4vGHHGzWfP9EwJtWy38HW9NFtLG9AZbYhWD8tinbZ01P07lxzuYgUZGE
FI42o8IfHHh886djmmqMzGUWOOfnk/uAoJ3rhcjQPWS+DcyY+iEBtKVh2fwyHaPNawxTdbUyHhj0
RxgfcJ8UcFIuQIT83Kz0DEwRNXUSpnvesEnICxaVqTs92C3dOXzISpyQQHzR7zlPMMSU14e/H8to
obU7pzlmHUwA7FQpmjG7B8sB6wWzIHcYd/uuDlmo/eC1u4L65T0kp3T5X5Dq3ltN7/HPRqKxIFXr
Y2IotmD4XXbVLja1WllYlCymPz/d1WShPhK06+2yzc8BjlIeFWVcAVxwZBu2wGG5i7HM8MZ2V/zT
KchnzahvcOweEGxnBiLYeiwIc1ehoGCHakqK8D6L1G6Yd4UEIPJ3mehMfmycyMEvxhWkltTg2trj
9Wx4v3p40lr53xbMEQ8XW6wRGBVmZ/swrI9Y12pzclm+LakLiH2pzOUEo/yQbm8TlpEuc2eicDCR
Ji6pDDlg8A5D8+B7NH7jDXp0YfQf+IZL/GyZdd/hTb4CpKHyNhZBURizDytPgVGsSxHtzYP1GJxM
E9XBeoeJP7FhonU8ER6fWrwRUz5RXDUD3D6rdA6jWcQLv4/tYh0r/0bHE9lH31wi69isXh8wbG94
LDGRpLk0k//0mrzSRnByPBpdtQjNabbsY9fOcy8cebhjtEYiUbGMhTcwUNUL+/BErO/Q9HMa0GUu
aSfRZuByZxTLuujsYQX5/HeH5GyBjd9oE3R5zffbl0MJ3MiCu2QjLh8fHRBwXEwM30uZXNO2Fhvp
MoONwtNzfNQmFpreZEKf732PICMIBfn7znPKTm7D44uTbIomCP4R8vuCidPrL00UVLKR+aZSFe59
rYNlTx/t3vJ/a3f2Clp1D3DfEAdKG4UXoC4rvOPavf5bqRX7BZz0UqxJREmtPeEHHnWbLntFFVnm
CTU+fuTEVCqHfnfIXCMnWX2ojhmz/c14b3uXhRmfw7nvEryCBhQV2uOYaDRPFzE7tWviOfHjNiAT
yGpF6mYKsjq/xrg/9fgVR9h+AOO60VK7ICG07gFrKodxMy/qiCZXTdfz1aw4UJJiGMBh9pSMAey5
9NyiMQPJNMI49WxtE6B/kUuRQ5cjrKNC3iygOKPu2+oGQO5CoU7iqR/I0E3ue/rlsqZlYdjUqcdQ
hL45iy/uIdjx9qg7abburFmzDfE9qN7+xj0DiQ5s+skOn5+gi5m5czjZn2Blm6kQb/VpiHvo/9JT
V+JYmQRXB9fnTYiMmdpkCJRBTkoMSS9W7GbRs74ULafNHG0UXbkVXF4lcj2tezEcvNEhDO5u5C71
Oa2XKEFatYfzvyW2qv4h0mEOjlS7w4Y2v/ck4tYqXuN2+ZSzygB9Fv8h5IkpAEXwKo2mxknvYMSg
9YD5hL0WV1mJLywhpegDJ+IHsOROFc33DiChtEQwKEsJk4VGIyZuqhoTZljBXNHIajs17V7c9zpY
/UVaNVa6S5Ihp2Th3pB6UBrPE5quER88y/qXNTwDOC215RIBaXAaSlIB+ayxGrzybZczzQKFJPuU
btA0iPe9kcx/vyoiaYJPvSUyBeyN+KvjSqwomKidEql5NHqu8rARYGhxq8qeGUKMlyUYTvjGRQBx
5Itc7xrknxrs6aT41MPYoAnyz15L0qnsNqN3pU88UdUf+lzmJJlwjGy92oVRR+UzJmLSv945XXNx
M6jGpx5xQc3wx2Ug1LIr09fJ2rF6sgpRMC8bK70Q5ucwZeLQ5T7JdOiQDGKEPTtBofQuELHsqmkz
R4qH/SOBHxO4YjBO2l9axAqub2alw0Yb9UxHypyNvlnngpbqF+0F8ebCs4iHb51YNbq5n4d0QsKI
sxwLqbgLFNjOPe6h+wtvGYeS72bh7ebT65CV8aYw5uhu0iOeRI+gIg3SUx423r98LzPpANZaa500
Kup+rxBFNUZD3jGKZPAejAbIdUQoMzuJwDO+QgEeUHReBWsYd40Ch5d9PsSLTv2S7SFFhd1e7UIx
Sn5/8Yet+LyBFp9pW1cCJqM/T9GMdyBvn+zy6+zYusnaD9m5kY4naUeQN2iEjD93OqFF3mpc7aup
KsX2vaR539cEIz4wD+JIH5eWq31bGRFszg3uFOmjsNb/KLX9mKo0ppF6+SfSdh9xV8/FF5T38FA0
Vq/mBmxHTPFwMJOFzmw/jLzHH6GseoT9TV6CU2td9r/7PABaHGbmhmfHotZpbFMBHd6uNzhKkQRm
FtEFfjUm428rlbAinBp67kuB7RnB79+YxrE0wl3B3PNrJwRXuO/NtU6O8KwixsiFslO6CQ79UTy/
cUUoA/3vKhAZE5IatWAbQ1XkUpBXxpTlZ1ULUyJc4aYBtsybHPZAurxmwrzcblAtF16vDqSYMWlU
INSxod0UKvntzteAF/kA1PT7hbDkJ2dZejpEOk5AqElGjZ/FaiZ4NG7HvHHqxUte7U1TU/CkXHJF
IjeN8Zz/Q1e4AuukkJRZ2vorqN0dpB5B4DXSYQdO9el1Yz194bwLdjvtbQI8XfViwJyK0F+/xCoy
ObIrd2NiQbrEKgU9BCd3LPm4vuWslmmWB3gWhSZEtmny86FWah1O97G8SoZ9o8+22rGvORDVG2+j
e7WyTJng5wZ5tJ/gsOYDJ4jL4nMYVG/nL0JdAs9tNiVbZbm1ABX/9Po+ko2os6sm3/ddBnWfDDBs
rGoUdiuJv03EknHRrBO24N2zSpIBcCECat6uXFe2WwnIaVcvUBVrIy0xKDfnHWat2RCkov42MD3m
J/cuMB4yCE0CaZstmhKAv6YEK1ypZ91EejEfEXdMtJwnVi91Wxzc6LOChc8c1o03v3IEnhLEvoMG
P3bGjab5NC5mvO4BCh/+0+Nwzn6sAQ19h8BztPVXwNMv+2HVWEaIDLyElcezytt3L1f3sNAQ5myh
g9iEQC7VUINXarpM1/fbHcCQ3RvEDDd6woCb9IKvdm0duSlEMEHnamGqb/gfVN/I8nHnHTW0GvhX
fpI+3iVeY7hTT88deVzJTgAxDptvApyaHZbKThQeSt21W5NZsaq5nQvSCCINg4EXkGJHNzdw43xh
HpskewNf/D9fFN3AWC21YrdUOxEU7vda3fczY6X8QEokNlV8BFvNWlrwB1pbptIeSzNiNzr6lMTX
amWpUbMzgdD4BCxRhuLNaAAUp43tQo8uwpqI/NF0Z7xapIisPxYaxPBomJES0fhuORar+89YJsPT
Ulzhq3BYcxN7XcMM9WbK8tC8B/HA7Os7OkxhzpiMCvHAA56V8y77Q0Az4wEiQmslmwafwTGPd7JR
oBttanjAkjboWvRmS5aDbkuYDnIg0wlnlxkFCuILZdNFYgN8jXFwVHoyI8pEkLtdg2Q+J8wJrbI2
8vdhuryvIPO7U1XTmPKa20Ucrw3lMpJukbXP/53U/xvZgdUDR+c1YisYFxU/DPI1OmRwtx9C4+BJ
nrAP2ePiRnamSSqO7n3p4IGMcfnEh9NniKjxNUCGG0asQsKvx92mc6olmNxrMjJ2GL0K2KT3Sx/F
1XxxJxngpfsrENNzxd1GcN1FeGFHauyrqTzGPAbkyH8fpjxoYlUDoDVDqbKeU7Mp0ezM/dA6NYQu
T34sYkiANE05zdozBJdR3CYGGXZfPYVXnCk9qSL5o5Mi/ttV965OckVwOrNDpbWi76/Vzugi5i6Y
s1rnAg4SadUtjI11QlStab5QemArfZGbCmmDQMpQXmjkAF7OqTDRyNcGNnqGSIDCxo932KwrRqMP
Puv+LQjlR9CMJs3Euq028aWb630VlsnBxVaveOlUsqpOKG7+sH4UMPyCyuCxLRjXMvMpaC5T9UGs
KSRga3g+ZtToktW761Wr6m5MRkTdW7VrhsLxVD6Y3UE5YgUCDtzHfKRoD9xMNm6icfjQky3ftxn/
GN/5Ts2OQP2F3JxnUXDPwAsRCndqdVypv0ndr2rSG5FvuS+C8oHhnJT7UQZ4Qlsb6BVOG067PK1O
UaNNG8UkL+V4XbtijNIDHOUl+4agoMWZhkMOdG0TnJH1vXT8imqFW7/sEHnVBi2CjUiLOU8+ilQk
Icv0cmrjVIVaM9LDT5SxsFkhkIQ2idkVxsfZKdAZI0BGRvkT6Vg1J1gpmeMpg22C9qvVJV4RG7H4
i1qdNVRQQJfASMy6W443Wy19p19IY8KedyhT+aQylhzoiQPBc3YOzSRo8cPpXlIZotPzU3U5o7kB
R6UKCkJ/hrq1NYaMwWe3u0V27+zbtlgzhTafw4cTkp8qOR8PMfhgQgIbb41RpUviuOP2l89+shLJ
btkAP+ICE7vSp/+kgg3OBErO3ZhmLkInQPs2Z/eYJRbRf32wbhflKFVGU/5R3oBXEqU4qRMxhzxH
DRLzT2JITp9wBv2BX1DyBJKUGRYMThjNVLL6n1CTxtsFoQZno7uSVQt5BMuSi7CII8C2YaghvtNv
9KsdIzrhOYv8OJJjedGKITETlLrF9y72L9Z9Z7zgKb9OZ7MGlFBHSxmMSj9fOK2eZG/hkH6u7U+N
9UNqAO3Op1Ps3n/8jTOWfYoHEGzVKeBSStnYtEpouUk6jB8tJaM5lTXWzhF1hnmQDoGK39PtQKRl
TCLqGRGSV+30ZBkTpx1UhrEhfa2bytOupL6D5TVVuCSNHK3l53ZsMe/TFKLoF66IFaQow1VephbH
2+Ek64HRauww9ddNvb8y9kX6GjJ8XHPA5/MBUewIwBO6fdIdQ/5nkjmUjP26ne60WWWQ9q2g4x0S
wjSo2sCq8oTF+8E8IG62ZpWxkwDQgsjRYhktZsJX5KbAnLi418MOoj4gcwWygfwgf51ceKhCPPLu
I3dA2MQ8HmiEGa6l911yKBnkbp7nUgyr2D0MgtxhKYsXIEDNd8ea62kKp1ptJgFVtfq4SiHf8xYk
5hZv89FSC+KfjXhZctVRPCSmMDLDLjDt9AvAa447qZO6cpai3LKlwqrf9k8u0VTFW+giGQuISVhE
5DV2+CpfZ7zpD370KgjPZjpkGHDzq59RaIosE5VgOC8uIkdyJNHz5IwQNrZdEgP9Taok0H2AgpwK
XkgGOpqt+06+PqAgsdTCnIyIzNgCNcA4K35VaH+5jSsbfBM7uyPuafPMkAiqW8eH04Vsgn/x4nAI
zeMVlDXJqgcYuAAttx21jiy2ZDUpr6sVn9wLGFFwm9KIVVE0BuSy2E08NNiHrrI36No6Vqio7Mrk
S2FSdHRQpx0Q19Sk07npAw/Q9W72q9hBUUCW8eG7xGJ4eSMVFOB59o1Tj0Iy8jccfvxwtcEYT8JJ
5akZL9vKYp0NNdbEalLDgxsOp/lij6qMSnHkLeEz7NbkdIdhT+rXjio8Zi7dBfy8jo814aRtuEWP
54rAP0CozFGfSAB9pbpZzihQ/qbF+G5IpT8dH+nmET6o+mlG2z3Ej8gQA+XfSpSevdJ44J/dE448
O5F/nE/l33EOH8zhoHG2ugeIhe50/W4DYscwV4eaqy2ZfWaD3eK4AKMZbi9bHdXjc5nMDcpRm1ck
yvqpq6pjy4lcrex3b8b3Pu6Tav0ERVDcZyVJ+Kec6C6BhtmxmzuyjDc0zArXCsT3NGNKRzjQFYuz
RRdlrSzRSxtrrhpog9jpw95nv2oT1FNLYcW9oBAFphUNgTtR6EA5AAMgd+a79hJB9SG92CC5WHR9
fMNG+vg4lB2XAMeoeAI6223WYAiNy6J4ReMAbZNvlJ0I4gigKb6O17Q4zpF/v4EcJOEQQ3HL3Ohz
9I9YWxgtDdtortEzuCqkL/7efKBcOprJ37AuxhlT6Ep+wroMoDCMh0bqjZ75ctVaC45ztQsEAX7G
VF93Qt/SAA1oclS013dLWDnxUlBdHUZDaI5Du3Z3IJ1Ii0ExD40fHBDjmIadsT6ytT4mHHmSaHu7
nlJDEOnav8mCq5PWy2oyCVKWHp0asjwZPoxGlgH9mfVdLb99GX8k+IBnsEvW5kDqyL0IFawazJ6h
WnDzlVKdk13Nw9TzuGm5jyR0AsIc47xKyo5t/omBEVT5TmLQRhb7BDSb9ZWFwG7arfFBGfTXa9Cq
OL66m26yfusy5Qu0AAQ6K5NCGmA3WffDhYqjnB/7pNsHhy5BrfabdNmMNI+5maTvOGWgzWjDeT36
/5pr9Pv8qlRqFT9KVReXdrxcl+9Cplp7UyGgPiEDl5srldrEyOOfmCn1Frq5Un16sv884e/pPxsd
ktvty6Hja9cJ8IZwKZP41yIAYGR20sq47u709cif8S37D3HRHgYnkz4c8cO48SNBYgUZxWdOiZOp
5FuBG0MA/kZXqk6y4sRZhWZO459N/g/78Mj3g09x/ZDoGS4SZmEMpB9HVcXZbaYGoI0W1oEtjl/7
dAUd6gZdYQsfTOAaeBvioupkP9u+vt038fiFAdsLcUp8XZvB0I662dBjqXbs0w/Yrr3Yua63QxuS
UeB4POZky0lTnYEkUyZYjT6PBAGIIyR7u35yHuisJSFLsCDD1kdHA1gJyiI7poVD8hcXC4RjXL4Z
3+slih21drgEnYjsgOYtsKZDPMPPPvF3Qx2MGQf6tRNNzuNLFc/xXAkMVlx9jSwMSHkt3xzCDuEv
erZZT94FZTQVuNbTxGEVcXrRhw+NNHjTV4aQjXOyS+g2zv+IGTeBJnYfWDOwjsoYfmpqOH6SUQ/P
06c+HPda+lg7RSERIoQMzYRwoFzBuv5Gd5fMysZG3dQohcz6RKcrmljb5WWL1+A4NT/ri7oAWM/i
aFwLWrvgXX/qW5Lxw/WophPxykaEviNNaT3pwDsLIRztyDvjlukgY4808z2BA5woifW3Vjkbi5nI
wTaA24q/TfvE+ht9a8lKfEMQ0oCmV8cKGLTs0/90s006vnX/NNdzMRPNx47EOPSurtIZwilbYJNi
SQ5HNz9q+3qO3DZy/eu8jhJ7YBC9LM4Ba7SIa+uBEMhNnTosd2KWMDNKxhmE96ck46wsp0AZVNal
+tg9wdDJCq6zCkoIhUNzeOq08/bqmPzYA/D5PPgQYkGX4TOg5DNP+eSoGuO4WIvo9Vf9QTX7ARGA
xVAgcYFvwrfiAAsGkGytrJHSgxgb1A9cDO1RsjxS1KmbPMuHWlYqWUs95GBk9mXdNGxmYJ0lsfsF
lfjfWN7oAP5y5HliQwpvhuJx2fRENNmgLfCvOL3zjP+Ehgfebs3AHRJdE/tejfj3rQx3Xs1g+EQZ
J2zsRye2dYXOnRsxVesoooB8i75Kray9/0mIUuxxbCsDaRZvWwu45P6pL6BNul8ntWIQIdfuZUbe
2Na28dhPr1nq/CloFoAUUnkB7xxbP56sG5r137oaq9SFyvf4R+znh+PzN0CK13yRT0uzttYc7jqS
4Db6jHHfWsNH6XR4RpppNnL9HwnlWBJTdWrI33RoyrPHjsrG5fpfYdxtmgLe3EjUOTj6QgUBsqcF
FCJxmYjRskQk0B1jfG5eY2iLnLpquZOGDGlGpaEn9RYduNXjUuoUG0+ggeZh1vEfInT7W/IPqg3z
h7PvJxecri0KDiTwM6CHIJk0XZbYgSQyzMWEXetHPAy4dsg1oCwfLqYshr/uXPAiXaYQwAiYGFiG
UkSnaysXBQP5XoZ+g4yKQLI4yYkWRxDJHBuvM4BTPKCKrfv2yeHL5rcInztKeJe57KG0zwVyvgMU
U4zuC/TdU6yjJ+T/urLyTCy+873dGZPOtK+VoRVj2xEGIPKKKoAffgsvOl7oyDf7EAtzQAfCNpo7
USxPRIAFfLMxozoCL7Ji1trqxQWExQm3vfL6hgj/Xccvqcy8Ib5apeWV66FsFrncq3pOaj1jJSTC
ewZifcZ9pXTE+pE5UHKOjGhf5E75Z7Qe+i+Jq3UYXpQEgXSBc4Mr211Iqz33rk2Q530PQYrTZ2Yg
B5Xo5mHOw3yTH25kjv9rq6BXMmPgzMIQafqmXQ6pBNPJODjojP4r23YR6s///aDV1pRlam9FBu08
S4nYbq1fe1epxKPn7r19yraiVOvHlRFNeIWuv+EU7aEZYe06IxcYFy3gQlqedmDUH88QNNfpMx6v
Ip43yxAFMMYMZwoHgcyhKpVcXDGvDxnLeKdpq/I8TRozM/hmj9osUi65I8vMWQBrXytmrOfhJHKO
juWbx0CfPbT/1o1tobg8TgwHdZSJmui975lC92WRJ3vkgZFbsI/It9JYd2z/nnU4VJUMfAa0zT+2
Z0gb1ZJFGAn2ZBs4YPBg6fer9ZMW2UcE9ugubphYxG4ZHxBCIAWnncHChly8VuOU9VgTxQlFQeOg
g9Jy1kyeyvhROGfEqkTHUV7HRBvpk9/e01Hff6kaDzEPMA+yUh8T+WiS/bCfSqDSZbYhM8Bp7EVb
/becyk0MHXYju21+H4KOZysUuqh58LEROIjpN/xO8iY/KuJHc4FVcg4WWRWNdhz21AFwZD8GIgix
GCEiivKSkzZzB7N2fFKEtQD3RL8pN8fCyXdDWXnCedvTczPhmmdSHcIqyscSc5uu4alMY6uzaAPa
guFA8Gtye0NYSk9WnwTQpbYteTXKd8URkqQOyQUXDWrRxE3aVL8k1UnqEf2zoJHbbFeyLkrtqPrG
kDAJ+bsjYTVLqyX356pAIHpAphQSlxfcbTVIkl72SA36LV+TQ1kduCJIc5Ryi2+0jJMod3wb5Gl5
8ltapo5sb0LJ3IidhHeUAYZvsyTSU6gx1qw7cg0N+mj4wnrInCE8Yhe3msxjDj1+jkmHnCQwCy3X
3q6izMk3YqNEzUvvbJHV2b6UVHFwqxuxTDqKi/yhFj3mPcHT5fvMbttihPX6eQ/LHhMPLqQLMByi
FpNdg2YV7zPEtNgfiUzvSnFYNKz6jM+opBAe6bIXtANQs05agM31NW3bvErdE6BXplqQYlPzqAX8
iV73owBSrhx3VP3Np4e6Zkcs0qL+rcTsVPxTxira4b3M+CKAW+ILlruKMjTL/h8t6O6lf/Vf8eKG
nqWgZKyRL3nBsKjHyyZRl5EUPqdAcF+GS4zTFnz5/YyiKOMJioWZhAx+RFRFuZXkf6aMJQXTjuTV
V0hnQ2yGxxdQoKnEn771nXB2cdRRqF84HrpMeQpSFBTCcE69DrCwVIzJpdkXOUAmxlZ6itRL5vNE
S11AO/0GNO2vvO0e4TituykcFhcBL1hNm2gIx94MdFJ6o2wp0MBjS1uibNBsy6EqIqhVgvAkvgdZ
iH+IhPPWoJCygeLPzbpZf9YmwllnMkX3l8oKtJgozwL/oH/Uynl27kUcRU4w8wZqc6KGL1MC6vrm
pmnZ9umI5Swg6Kdvv1A2K+6F/nhfpO6SUVnZk9ZM989HInCB7fYcfBKDy2KFQEqLCCym8yzrj/FF
J8KV7aLbh6MQI8Q6CPWSelrJIarzGkjSbEuYrfkrmZY+PF4RWa1Pf0qShjzHkxrO3Ksnr3s/INAH
NvxszNrJQDJ5Tn/eCbWSLJKQNMS2BTFt18YTOLRctHq9SaiMW+2Bl2NS7S0WUoulERL8LqGQ58fN
ZgceBWSL19a0PzwEa+9y5uOBfvkMeZ3hHxzx85vFv0EBUOV4p5hsAwjXDzjImpy5qKbYpR+mIP+T
UOXQI5SZXinOCnrJgEyR4dFXMfLcLknmwUz6frGAEamhYAjQp1C7ujDrcJj03rDpV+GXSDBluX/D
vRz6B50c3P2S7DU7bzoKXxiX3fJN99zhPnh8GM6w5VuIiFrEvaqKZkShkZaC692iL8fN9Ab9MgaM
wE9DJgeK/ZffJr3QQskHoV+apbLB513DAGVuf2p4j9Br4iJrzTauh1lJGiS+giqJHw2feHyVlWOu
AB63Ddk9O9yTAC294tD7hLBLlNJcJrkY5IV59GS7HfMMp2hpYuCFjXAKHoyDwOhFrKFx/epLs4jv
Xkq5aO4wDnASUiai6b95f4fbxorZcw6B+W9pF1nQ0W/Pl7AQWqN+SP25pHKCycNPArPl521ZVAG6
hvIkQxa/7BZiqfMR1pu2R5WIhFzdZNOXvDvp9w1fZ0WpR2HAK0xUqTwwkPk5WS0EpX7/khyjLYqD
jSm9YtM0HoyTiL5xRGSa7n/SRGeiN5oPaW52cfkAl1C9yAbZZAjWjdoGQfGHFxW8TQfE5xeaXt6J
yJroOo0HCKn5o+Kysii/MtDEOfStExTYxxUNdNEgsZFPDdEZy8n8YHqOrNUUUfkpYqpiLomzObms
cQ6j9ylVLczgcarzKgdKOeSrS3reZkflvQ1YV5r9o12O01QD+9qkudHcRjNF2m9Dj9hbAnhryULK
BLdri1ozYCQgY8IsVTODm72VntgUjidVzFMv8RwNlyjH/htUl9kuiua1E9rj8r0eTMGR/75IySDx
M6S194KE2IeXqP0OjbQ36GEZa+UAJkJSanDE0zgnENrgW80OM4i7VuRx38EW1wRR0CvYJJdUbtky
ku0zHxcBoZpdkJMNVw7CYTmng0EYnRR5A/Qwcn3tPpqj0aVPKuDVVpecGCLaicVBmfbsgLMbc1po
GQ1gui5+OdTo//UJ4o4Favg1n3nz7H+TnW9FZ0A34iOKKnGjprYFuU5nnTlROXrUU9d3J8+VkeM7
sE5S7A2rgNZEg+qzdrP7t3L46BF9gLOd8T3KrzQYjTjbyyUn0WgP/7KNIKnJNzfN8CLQRCyfZXE+
Dm6Xm1N+ktQZWszKH9EhIfBvGMElL6W+MGe0wg9ENpxtI9kChk33V9mGFqpcJx+0jf5mvqRJswPw
xkiGKw6VSRmnnqKe0V+3lehcIDLBU4nRwWV+dIKFML4uDA0sQ5LO5Cz0ckyI7vofg/ryE1nvZWvw
QA2C9BITdYXhtUTjelo47PJ63jBzc+Fe5osCeNJoCWreHGCLXgUxyV469IcNhbnE/KwKU2mIAvgg
cL9M8W7F1o4kiYCzSwmpSfFABJ8AaO/cISSr9WGjGN9PmTAfzLhJXi02aFW2EwIu1JHs63oUr3WQ
tW1/9VGBdpioclUpQtY/t3JmikkIf22vJGbVSTHKSJvxUakmOLRVWThZNUn+IOboikYeuc/1oZ9m
Zf2duQ3pNdmx2zhpM26l1uc5gMx+C9ps+ra15E0A4UQDhomgxZ3fEuPlbVZqySjD1Rj937RflL9q
kkvJVZ06elHYjJVNSlURbuWouEP6W/jgj0rx0+4rsDDtOhaUeVQMVYin0jgxGJdbH8Pt6YSWBrXj
8HvW+Ai/eqfxs36lN+1+a78BH1EZYpDtFRtd6GTmpT+G5apfvQQUTZ83Ayop3UPCrz5V22vHIVtS
SyZtqhDop8BlzAqzPqIQ6rNlX/zZz965yvHKVuUlYAkosV5L0z5w3zAnqQPGAJGjQ+rE7mOOPOmz
Bhb3xmoYQs9Ro/UxDuqyYALsY5WgqMkdwTlCzvMNpGExvZUA/cn1PCIdhJSVlvJWKCwQBaAtoEDd
FA2NilOWQS94V3puQKzfrBdmqvtztyCGb9d49LRy0OSLagC4D5hzmZkTw8155dJ0MtGvAl4veGOW
NtI6/+QIykRANFQn0KLWyfLFQ1CaRL6mIBsO22GsfKrIKYAazfBEijVk5LyFIh6s5wErbfqsUQWz
3xuhYv4EJKnaSLPsCo4uZdzxWt+evlVN8rzgpqyP9Tk2yR3y4din427IL6U4wNPjN0PZ3JXOYV/K
JnJKoPre8vfc3wFgo90zoiCdJSbusNxi0FJAIwkQ3OY8FNkTHqd6XmjSaciB10ZxpVu0X1dinf4l
0C4h656foLMJSwvhhp2jZH8GIRDwZXLWYAOO8a9E+YkO2YODf7tfZi3F5mQ/WO19UXjnrP6HgrZx
Isx4OZRCrg3HqknhaoDwBlYWFjsoKltzS4CwaqLstUKLsuC2BxGh/EtHIAutgdsVzAXhgtmo/agF
y3GS814N1IoOltLlo8awu9hJ6oIbMlSF71kgN/BJB04dWvancBwYwgYilyHclFWF9/z0hQ6wrcye
+3KbQgdnGJ0YEsnyMsMjm65FtzY3y3cB2t9BDVtd1KTV9JHTMtbgQ9mJRqlkqj935C5lDDsFR3P+
MccPbPBdWH1CCKGXV1kHtfv/wAP4WmlmcpmOPQuRA2fAku8Bc54JzJwpjg93UlhOkWae+gOaVp27
EiFFwyKSb7aa9qVge2ncQSBBVNxDJtxL5X9mt6pHDV8ekeXZWzr+PMonnPYbNdpAsXo1K8vlSb6H
0BIp3cP62j0BO0TJ3mAIDQ+dpYxBPUxeQG3pcqL9wb2Jpns3DLxWW4askIitBgEqD0HOiNFz30pX
n8+r0muLOg36J4+k0r3lOix1KF6rSws/RGVTTB24zIxh3n7HtIGk5fRTr+uJ5auOvz1HXtuyDYr1
aTzCOw0+mp4qCrA88PUoQszwxvuYC+pFc7AMDPULinNSkPB3TVvxpC2cLPHtaNeShz4yCYkProWl
5rJsibfhQn6WeLwbZYjlYYiEbxyu4Ei3gAf0RBTs03L4P70Eu4ioV64RDOWHPWsqxqLXRUyo4c1R
pQWL9BFZPSKGkbTAtPr6Ty23SWzGQv3+YUOTAsCw11UgDOGWXRhhbk/S3YF8dtPM9S+Vf40vop4X
er54igPPE/5bvH5jGSqXOZoK+AsmGFUpgtlNfdrdQAVQLezBnl/wD17C0A/k3JkIL5WaXUHADVpM
zPB/5G5WWUkMFSfK2iHCJ8gB47Q7GHoxmwNl6BHSc6Jf1n/2W7/DC9WuNyknSvsYjIDQi8dOFq68
AKPiMJYeUF/XCqLH6k1tvkPRW131Goi30o6K26AUFaxzvvuMnX1bbCMQ0u+Z4v7RErhKnRVjnuIK
Eiupx53l9Hhj8tgsEkRmQDMuXjLkZJI5PpLqN8Wne6W4uW7gWF4YigdJNZpHHMSODudlGrHzjNcA
vJ/qj+uZxGP31F3690nITKJiT8PAiUN54XQFA5enj4ltQ30AXi85/6GMcsGbnQ4uKog1Eqf7527S
0k5N6yC6k48YKB/L05YC7V5TVf+fm8SS0tf4gciPqLgN4BYGPX74sXn9B2WJNdMkaGxYNK9Bfp7i
tNrsHKypC7wRf45PrnrqV0/u5ckAYS46TM75HfiT/8yKIeXJ+2kjr/hYiIC1RLuQ89K1nm/BMp5w
NPpAjfdA5/mDcpHf8KPtI1hYZ8eZHm85/cS1/VgHwdhwluB8yTLayH9q+HU8ngkvJ8Pwrtbm5wAe
Ug+W0M5ioRq9iq7Zh5EzRqxPyffYUPTZ6jt6YKeymgHt/EJtc1OlB1csa6lyi0gS+d1Z4Z++mktX
vxVEsrs90W06JKWMM6hyKfeW341GDkfIO5lTpt1qJsm30s1w352AMsHy47LDD7rgZ/wEfHjGBf0N
sUAurHtgzuhfoVWQdfC4d2fzCQ95IEpUtbvVMsO85PLlvXCGM4uchwMdRyDQDN2dgmcqZWJXjFPL
xMP62QVn42PIWIGFOvG6SYJ85jkmIptFl/SveV08OV5IgIS3ECiBF2k6Q6J9exVQ9ouXFxk4YP30
kFMTG7bbYpkepLhXv0vucvf+HX5LRT1mByFMJrRT2pcBNwzEyjntkVc7s33RCieeEIvn4tp/rv2k
exVGXfumDJSuky2CRAehwM+3+oxlZyXQ39fDZZokQf2ARoUpSi2zc33sW6L58Jah6pYiMl7o2hXt
+3akOCxTH32SB2iyA5/k70xnuCKFKrAeTzFEhfI6a/mt8++/5I8+Ajr5afewoFE/isrzwlptu7+J
f37kvPOWQUqSG6xNdiEB6ZAdYbvP/e3GAhnx5BgI56JlqpofPdaMSyNA/qlh6iam1ug2owdDfxSw
wOGJDItogvAofFFjxSbzyJGMeL+1pV5KiWpltydF/FQsWWCVfYq0uetBvVyjgcg4dxRQ8nfN6jbX
s0NSAEg6vLHUurbRz+QihrxnVnCOLXpB9crMxY3vPujJawd/3UcJXXsmtXWB1ZsrngZBycXhkmek
7LauP+PBfD+sdJpzX2tkihp4OPB62EKfqc7muG2lRrKSpHOnJcCinJDr87fGuJ70SgCUoHAqtDJe
FZbbyEheLoH7WJ4I0J4+k4KimhxqC/gWfRIpvHu982H+Y/8VSqksTUFcM9mi+YlDoXPpFV7zB4Wn
++GWj46ccuXseSWAtj8H0QOcaJiR8LMCpzATTS9tkDl77FHWA3E44p21JoOkv/g5L6ZQubVZT2Ug
6/mHmkSxsjCmHky3IQ+BCiYzYs5DpFmkv5rE4gzYfFt0gX4Ql34G6IwmChkspGTqXpEeY64CySFk
CdOEIeB8UB0hhK8LWVgDnaMdMCRcNtrkWz/Krwtfk4OWN/2HFGfuJkVJWBgKQ4MP+v2WEKFEZTSc
+yWWOWVT81I0hkpUTvxj4FxQA6E3G/sxsJVCfIH3ga/kebr93YPVx88SojQH4Obzu/lqbo993HEW
6jll9oPps/N+JFCKcVVw1/BdXzX7i0Lvd05ZIIBhPct/OjUmpPD3HHhFsxwD1XhJIAUdHdlmEIoO
j06AMSptvYVEoUB+ox00U1iMtPqAAtdQKBKKWAK5Tl/0r5s9lMp4T+vmCqIIUtZdnv/SRTXdbqYu
SY3lcWV2JbU/bCEHKED4uVNbpRbiati+m/4IjaG610yftttQuT9lLYtl5sN0fPHVxTMwPyryB80R
kx3aI1BQ3xMCjVxce6NRsFZ3lmowyKN2JYB8HCnplq/86AYx25tRR2CV687KHvhkPBjzIB8f3otR
wO2YfsziCSdO8JKFSxdYGZYr+Nq/XoAu0LpLmyV7hnixLg3tdqrE+ge04fxGkjvqb2vEtm2260wI
bZuJCAmAmJEm+y1aDAfYn9MSUifqzkUHgalyczdBoUCkZSGrDNnRaOkOe5t6pi2J9G6VwpiWxgD2
BGpl+1x3npYSMLmxEZEEPi50yFs2bEFwjowyEUAe8RGT7I/s/RvLrDIzG4RJJOS8gX05EwuqBGfh
tUOioW6CuPTeKP4c0mjYM1gjvefp+WHY1KJn86Ns6kutHb9wa/ohZejZRpyietvbKjT6bX3qX+Ee
tuImrYNZH5BTywsobpoqnguCBhqWNMD1myylI5/Rz0EKZskNOVQUXwWc5zMyz5glZGi8M5QwBPVj
yUmR6o6F4FqJ05YtvbTfgiKWAXA5TasBFAYi8tx3JVQoN455HqWrAREgMd6Kr9sSBITtp3cjx5GS
+XHvRFdzXwIZhq8xDNGGfMEUtw1ZKttAvETeB45M1is2r6b01AHhmvDPQspJSrjwTBvAlNNU4FFJ
12lsEC4r9zmBxddsB+4QghZoY21g2U7G4B/GLhUKlvKmkYWP4yHtOviq4c8CCqgrhKCLN9uNY4eb
hAOyMrzVzbd+3GfkirR7oJiKLFwl9vz0rOgNXTIr4Kz+1GVlSK+b0J6SeisUwd3CFacqjlodi1Jz
rKmTXcepmHkpuBB9b1ZSCKi8pMwiCXx0w846rTk9cgj77OK08+wF29rhMxK6zpAChapHPzYyS7gO
DJElhwoyY8t+p17R7q4AkhLL0StSx442svK6Wy9XKZSwXfMzhpEhzQIDjeI6eLkrZ8j7wcLNP3I1
QsGlaSNK5LaSqITiYWW2AOURdEOMgDMe0vhfj032Bhz3l72iFytQRF2HrMHYl5Yv1hS7jShIKSLd
NcIDd87LWjuy0noGBNsWAI4yt1yN993NyxI0sJbu7W7XcrWXiKI7iNRmYWUFFHWiwrj4RUvN+W1d
Z+AEXC2MZVL/sU9PrVYVDFQkj0NAonDTYzE95Ii41cdpLp8hGttuznySabrXOiw2lV+f/JKqmiBq
eCnU1XfN1nZAa3H5V4hIApbJpQmmzhry6ZxRuxJvCa3qJCziAWRdYjWymh5yR4MqtDNKx31HFilT
fj42hkJgL1jIEPIAE29Xi0xM17yWHdC0Y9PJBQXKqq6sthmI57kvzsXQ4WCJR/+41A5obFeAQGRv
mIWW24XF6+51ogYGbjEqstlnMtcFsL5Umhlu1ozgSA6KphzHkgBRC6Vckj5rYbX1Mj6VV+yP0jBl
24EWkSeOI9oKqjwQJYrdKigRbf/Hw6KRvWXq4wIxyJQwvM7UdBLzOoaMwais8xAWCCgxmYrF9pnb
87EY5NeGmEZtnbB3Bg0/G6hEnu+6ZzqyCXDmor82jkkaNjK50nsDHA2Oi5lM9JcHwCkiNu+8TbS7
zKRhQJqF4lIGJ2+NKZkthTregEywCp6CXf9aS8TzCwz5KN0novc441zI7YExcmWaUWcs8o6aXq+j
dKtfgBQ/pi+H78VyE9OCev7J4zj5LnGHqW/Ypp5wRtI0LEFStTDMmd326p/+IaiJ+LmWW5GqPVqE
WwFUk6iwEracw7P6RBt87wip82ASD4I9l80xhrouHSgtrOjBvfklScwShdxtI9NaNlnKjJ3vRhEB
avKsVY9KjnMu7fGEQc18AGC8zpGCH3yhdOStnX3brqp/kXmTYERoujNjloxLseP/NuNIPCDO3edN
h16Q0YF8dO2lPaWf65Q09YkTmqFNR5Ri3cS3g+QO/hRgwyq63iPweAVZp1I5rQ8BzYtT/GXMQe2m
aTV4QCXWkHZa0Ggjp1tkfGFvc6luNVeBKs0Ou5+7utIvklu48NktnkZ6F2k3AtUOzFfZ+vir6mQ+
YvJ2Gpxx/3kP94QGAMmMQazWh/cYiuJtfhvllFLQPV6cbnkje/m+6yn/0UzBjVvl06Jmh8A07HAk
+R3A+I6ya6Fqb56SqSIGA+6qyr/qdysuAa4E53JzkHggpd2EXgUJlBR+83S0MW1xK55FZ/vB/hd5
XC8bz+itkVAwoZEHA8AZ+NWQDXtiMIjNvQwbDkn+LuUJ7HA2psyoHR15itvGI+fMTx12PV4738fs
xaGRhHnYpVkmNJ1KwPA27KD3TRnfbHUNyGvnVikJx7RJwvbpCgg9h9n+MqZBDqS+OiEeLvH4w95F
2hKCvtOMVvox70eu54Yn1jBGcgy3u7XpyDJj5jKjF4CeNu99P/Yk3+Ig2NDD4iojEUJ70Uzw/lp2
xGNoK831I8r+6R8vEXeL2AlP31cUHBtUosjJVFZ+x4c+rFIYxVuCBBG17yEDbGKcrNzSIjrgvnyK
62xp4AAx7xpO/zel1fG9PixwNpjLVgk3kFQMrFR/7fTsfF/GpcyW9bMy3HrWBve5OvS+yvk5Atdq
NRIPbR5nwOFihQaIrSE6rxkBIvKM096GPuZnwiC6Y0d0lO+WstXhjqBJgckbvLYpzvhWxP5gs/e0
EsKSHTQ8Z7dFowX/tav+9c1kyJgzrJCzKzPqlN9QzNe2ihES2zPmUKd1JweHSU/cqwFsHUAHXGNl
WIuZE/p/gZw3KzNCngFKgMAYcdGEICbOuOycLSnTehkT9jBrzTt7cEyP1EdRrGnwQql9JQ0cjnE4
dw93JqJiw8bcb7b/PPZsswADgx04xbaF31DgRZXe56fwapSjQ9b40BO1+ay+iC2dEHeE6vstCmdH
KclztgqLwUcrdbQjg8/uvkQI+XsHwdQYTxyKIOSEklJ16JA2ufnKx3LXi+NTJ9Xs6RswiilA5gPg
GDReMlF7tZebk1GimTtKr32wOvhc7NKxMFliq1uNCTvLwyN6qV7tLaV2dOOrxWNnhhEEUucyWe+i
rxG/WPSTmZ1+JDJgT/yL9FaCuLV6NJQtOfiazth9S5/wSZlYoQYIvOWhVRxoT+Viq+0l8PmC1lY9
Iqy+hZwjW1tS7GzgjU1cvzZfMQhopHvd074+LXi9juQgpTl+HnohBIMXOqy5vQtmehUd7YOcT46Q
m3B8HmERVW7cSTnHj+cvLpEld0D6O3Llp4kMfhG/RhDidiI51R9ZW4vj6yCH6FBJxEpn5wxzrxAa
7PsW/LOo6fgNbupS02fgwGJwS+KmOePvc2JfP/e91ZcnLqC9vGsBMO95eow5Zg3wetGefCr+G/OL
LGpVvLR/uZSWf1+QmCJuQ1JHqyyHeKpowSQEz2kpqGRKVbxag2Lkmnqse8dlafrAgNsJ1W0zDktj
GoDYYPF94pi0MvR2Y+m8h8pWAr66iT+6dt94wbVCemp9B86RK/LDw7hy/dTtzLfkOmbMoiCuWnyH
kYfBtHOnvz9d/ihPWZcx/XTDULIhTvCBQIt4UaZ2ypj93XxVGMzrpj3IWRoAfJ1GxEvuUyJ3OLbj
30gAnSNlqevFQ0wCePXb1/18ck2YuUieaXV6AGUxH4uPfG5CzF/bSswTUEhEsrlUDk7BHXtqE5PR
5iP/Qu2+fHGyv1EV93kJ/V6f25QhfgIPtQ+zAGfwqb4dXlElS4WTKPpEtArp3OSXzoTCU6C0zU8p
yEIjlgoW9StiTI4DK+uumTAW961DLoUatYApT4vUd4yQASgO+vUZzdYpnGfdGLonEuzQQMpIyaPb
Ur/Fnt0beJ3fC80SFsH6XRjZGMjuudi1U1Xi6jz1J1S92dfcwf+E6DGVOZTVbOO6J4Nekro2oRSu
sAWQHxTnWB1l5mtNu7kaeboPdAa/KluOt6Z86UF/LFhzQfKod4+8qFfrtGytuN5/+qz5ruwbQHHS
m1FhaUhzV+i/Na/+TSv6F8RnvEjJXIEobD2PAxHtQAl0O9x2kIJfJkXsyItMWaGVogS52i8XpM/K
qgzfpqJ4CEhDcZ52kZIP0by3ULmi6zohw5QG97VXFKKbJp4hFyYyGnu9xi7APgb1l5wE0P/64CQv
Xv54cyGlW0vLTRGxu+sUAuXee8LBc6zPh6Yw2EL6CXoytLHZG5SiYUDR0hcv1dvbCvJZTmba6Q6g
NUbhS0bneVpcllTxoWxdQiPDCOgA7ZaPMplRir/JYmfSNOPR0a05piuwuDsPm/bQzCF3hpzbKvXO
TfqvdbW+3giqGhdvtJFYCTcQOhbqm93gUHCL6an4QXgD8P/z3c1U1O4Fb/8dO/DIYergADkDLFPc
btqkhMIFVaaCs6rC6S/mjp1JuVjxdIjSDvBPtB0O6snrn4UwnSDYMC4QEcPLK6kcpzM+crkgvYgA
VvUUoIN7Qp66tVqyn3nVsCb/HPq+RcdU8l8sc8vcAztWCRqR7dkfOdBtolip8BPSD6g4e6uswG4t
pC/lJjAJ/Kuj8DvT7NvOpDnTJ+5isBFjSL6ZsmfKCau2HRoVhOW57+bA4Pm6MiNP+mMT6pXjtHEC
G1fJ7eut5/gpAN2Ca0eCSPr+eMi/EshhgYceM3cQyYS3fwLU/dt4829ZpfxMhy4Surk8wZQTs2pk
ZiACXGS09QAvNFKeK8AH5Se7xtcSK6cuwktR889VT9Wt9d/x2TQibIJjmTPyY/A4KPbmT4mJc7Lj
zTKsDcKb5tlPpT7deqcyEMV8cPQs2aMihIDgY7V6NxzM3UhJ/AcWUWtpPfCPLPqmiIWSZl3UQwzJ
ku1jZN+chRARwo6WKDBfRQNZWH36C4+O4sXrC+wegFAxCxm8Eg8P5c/bpS5H4C9ecVA12zF7/887
ct/GYE6bdbf/i6gZIAD4GQQ7JEi5qQcPIJdCxXGahiOWNs9E+Pfb8NaP2VcoU48ZKrjMgAGIRLlu
KcVQbnDls7Mlrvk1p4YKNd7YIsR3A7Up2XeNihTob9WJmpORwZALYHjgDebswpIgexfBHJggvbI3
vWmul6ksJnnWTDe89ZfJ1vMCHh9aIV98FdbZWEBdbn3fT/1kO3JMLdZjGuZSm7al71GdQXmN1/lU
8div2NZ/ZzytsxRPAaZ7moc4mDrclIgmvWp/vd3Zov+wauQmgcmAmOaFXI+lb8cdIeRUjBOPUAbP
UB+CAJYM6i4lAdBW4qvsQL/xfhLXImzQxFmJLcuDzS0miUsCBOkGMEXNme91Yv9KfJ+JK3YEAIoi
czmWLqV1ySP2cjrISKPL6Z+An0dRPXQoUciK0gasys0Y4pMKWHpmn23ZO3VKD3ft6dOfWDTw6VHm
jeTqR9eHeqYHnemfiHQyjvz9u52m7CtXu5R8D68wr5DzEgtaNx78tIGp853r2gyTRV5b/6nPOWgZ
i2Tr/oeRNROYBDvCJ5LvDHWt11cxzjAO2xK3xaxXyy/qCb25+pFLaXujDxedLZ7smw6MSO9X9N32
AWFkcNTRdcGxLzqMxWpJ1yggpm0/HyQuDQ+wPeMzWWih6t6z2VKOUffmd2pXKL8283LB7MDzRFlS
3n2aumumBNrOoSPuepxrsCVARTtG7ciU9rLSjr3qub1xIZhTUjY9tHIClRfND6O3LqaeChc+g2eK
nLfmtJci42Mw8eUZPoCIXXNm8iOC6P7g8K7xYRz6+7gcwomxnuykGsZbSwq7unqiVu0lwL2tOaFr
P2sPdYB+0zYRNuyDZBN9TsjLV9KQREYXpa6obd7SrJL9heIunyJScxkcIMPBIP6gxtzWX5jDjYWH
foI5HFnMHwyf/jGLLObuUQzwUc13H3OpygtF2MvaOvf17yUIIcMlWbh14eze06KbO6pQeHWwMeew
8qhPYk7VtFhe3kI+mmBqDCvrFQvDZrnIrMdKJnRCoeqUtwJzcgGk638IM3v2iUihiJ6MC7Ofar53
S4J96wUbfXLC68Ng9yFZc+Ns1ynqMg66vBPdGEwwR/Qa0n5C8wJ8hrLgTMT22PirAYIzl7CsQwjd
FaM+lJAgSvobfHpQu38b1xgjcmSNECbBhr8velKJqZtuHKP8F+n4Y52NOHZmHyVlVDGlbet8n+Ag
k7C54B57GlPKjd16+5tt2C9B7WV/mtjLhhRgMQPkCsPtQROioKFxQiYfFNuRDLf7Tr3heS2UUAss
3xSifENAxmS6M3L244kjVHEPYJygxCX/deDxCnSPgdAwaglmuFt3JPBWeFIeyc9EHV96/0iFD+v0
w5mgzJOAuIF/O2Fz9h0Wy9nwiKj1Wr85nPecyFbFhJyE6zCYPyXPX1DXibe1gnAiBKamLgCRbi/m
X0K3thhA1zZvQkISYp7tzll2+l/A0C7hgWQ11n6UUCjjG3jQEe//mHm9GCszB8I9ee9xJhIXq/gk
Xs+m+fDNMTi71WJk8icbE3pxp7QGsdBIUVubp7jSVB+6V7D+w/MSWYsBYRv9usV3otYbBP+Rx5PX
zg2kP7ApRyMXsNK6beBwmqh51BLSVXM/sJB2jyM8tJOEsitJcMFwFUXFw1POdzOmfUmn0jQ1NoOU
dHUUfXtqpTcBV21twtGlWqo6GukoIXU2u8FH3x1oXOrMqWVG3oyZ6vQldV+A0q/F6niWfrkgn8ct
WkvvvNjAUJx7DLzf6m0xAYu7dRht5xXuIeNDAKF7podCmCp1+Vv2Hpp94DDehWqyuE/5QG7E0pbU
F5DGH7JaMH3/VtsqYqcpjpdNe0cdu7YkWf/6gvTynP8kWTlKd6Y/4XStfC06r7+Z1M/ZxxJtE1t/
vQ19F3CiFss4Rdmb5xsHJ9HqxT2xkjya38/4E4lsljNzreDVhFpgCvcFyyR6P2oi+800OA6dBe7o
uSShEakGvuupl74V2lBTz5X1vRM+a0WqjoD4zA7vHmYsAW1mRUZ/467x8ssqCuVf+lVTuZY2et4M
pLPc57CkYUa1bDLjMfmZ2HDS2zTDdBN8uhoY/hquTOnrZiVPXnRYyVhui9ricM/6k5QxnaWrueoD
IAFXzEtvfHqiijNwwflXCUcI0J8SB4VuxI9ru3KR2BAIvcw3OuHTlGN+bYSkdm8U8mT9HPd6/dgF
lsKKqr6G3gZwdoknN+zHVN0diqahQVKELDhl/qgvidWLD8ZP6GjZaufjmhsAiArFMVEdLsLnDDNu
2p/KdNyqqBL/SpJupiAroiN+OVYnfen56mZll7S4rcemKSpAKYNMZ3igqSNWf255/7dhbUvUhDiq
lXpEdsVc0N+YShplDsUVMIIiCUI3Ul6/mjNiamiK+aHqj4yo2zx/MnJYVHlRSMaRUwJyWVc9xOgD
8W6zfbBLAvurpKrElXL7iZLyZw+65UGuiOb7ZgpxlubZoVUjm/6AM/Rs/epcXEUAaDc37e+Dildg
vKUEtK4dWxTk6/S5jgPwo9QSW2eIS4dCy+bAX/ydP3ht4ryyro1AVkA9oRQlMkxJIyhojxq/f9IJ
gZazW4BAUhLMGYr+v4dLbeuzOgJZZCzRKiehLl7UuCp3Y2t8A4Yet9fvTTwvXgDjUNJuz4QzjBt+
rDNwyDdFoa+K3JXy1djzsBWYTg1sZhnoEJvA6cuQ+5dyeIua6eg3jYiuQGjbTr9pITzAfOE8G6lw
bGYJqos//z5jHPdHfr9xGzdwuNgjRkZ7A4hQR7xraSbhLNFPrAUTvIICa0itYzZpx1GInvyBcgbS
nDAe7ou8foYPoIO+S2eHauomNyUl1kVYFSGVJTbbyWpmNRhkt1qpLqctlxM/vCeFOuVE1Kp4KCXu
LKkdV44GtXUeUFZfcdA8aBxJCTnUP/Am/2o//i10U04UETfIxhoD2AxIrBbSJ3n4S2MGGU9Nw5f6
DfTLejtd+vHGA+G1fENz7DsU8np5zcOKwgzkYqd3H6ONEN+9MSvrpEmBQj3tMsNt5RVC7+uV6kgO
lMcDUf4WT4j0sSI1bmhWKSCfAiAdHMOLZAGKDaaXz6IvBiU19vyfG+59DKFF8Km+DNOZdZK0q7y6
UUnzXWZMoZKllJQhOauc4HrPWO1Lqqn1dPRzRWbV7dHkpSWVOxXLjDSNjeBAoScMT67KDZwBnI/3
x5VEj9mRpS/w3O3o3AtECUW8kmZ35pvxW8eXzm8k8QgF58PaX8g0DaUPqjV16uUGMLcKewneBfdp
BYFF7cgL42Gmb1FUsaD3DWI3irAIwIe3gAVp5XbDue5Ac5YKQfO6She2Tgz6RBdldub0g05fvLrF
PRhUu28vGdB3Eq9DOdZYIV7wahVyUvTCqRKGk4jC40z8wx1YvK44S5SEMaWKQhFbsFH/2uwoVmUM
cKDY6MNl1Ylrc38aX6qM6MeSQz66j+gSrZdQVY7fOuKbOEtQaUyCsEwqck0m+rm0HGLdLeveF5Oc
dQeMn2vLxF5nfVbQnul8irpLjf6muGNxL/ay3G1OnrBu7NVa8OrBI71su6Ijbt1omc13gXwukF12
c5tA1imYbUStT4r0+GpZHuqAXGtGBdxR/6rR0qU5Mq0JVPqim+mK+9aL5Rw8WW0Oy7INx+kKzpNo
+gqTJPlSuH54L2txt8Xlt3ZYo6nnaLoFgJ1zRFaGvPaAhr9e3Sfn8Q9hnYuDceJWUun8/X0wMTde
KmI6LBAgRKM3Ij09IxAYMAX+jEBPZRej4lpczPGAJ+2svVVqyquYlRuE42E+gDt0y2Oy/HeKphKI
jj0awQgrZtr1xAgLhbTLhZrEQb46ObEjBuEJAokTIjT483+GdAOC+nwL29sgq4YePtnEzgiBmxyi
9B1O8KSnbLJ8axfcql6V413kVIGxeyhNjoI9VIwvZ7MAslB3oijp/AEtYx7KpnaPETKV5ZcPMTJe
s3/TFd8byxql6BXgGiV7cORS0xrgsh9twxIKvHakrAvgrumU7tB0xR/ut6Jdfjgb9Um8Xcb7KQfM
mOrff4dsJvVhfuMsKyph1EL0x6PPMKKBPyrdjJukeJH52n4yLMQbgTRG2RQ2/eFY8ZpfoxPqcPc/
G8HnKemaK3+DRkylt79eilyXczUGow8LzwgidespScPpHSdorkR4c3Kuj5MNRQt6/tqR2rhUPBW9
FvCW0fcmp56JtbBTweHw4tuMZUsUbJLjr+STj6G5qr/i5hOUhwKW8a7sr7n5Ryctyi7UEq+k99BA
8P6pTzrCD4eWAsJaIqvPB64Ug408wk4hOcmbJwkUlfhVxrFB/knR4F0oz1CtzStDYpmZ7yV3Ak63
WDL8F+7Jzwjo+MVZkN51IlDLGQx9rhY2cVoE2eC6bj+4iCmKHjHwA7Yye5y0q5RT2GmCxflip/OJ
1NIjBOQHZHb4V3DF5wzsqPxhsQpWpfCQvKHtlM+M6QVRTvcKBL0mBIm91ioPuJMFE6mPjAc+TtvL
U7JnkPVv6UMi3q4ye1Ol2XAQZyrzuVhvRupsQlTJV5VuQ2ndIVxocVhw8vR/BNpdsqdHBvAiRHgh
JzAY3KIzpyjBHyjep22soXkfLrxgcohrQDNy5hEtrAkcIvi45O0Q17NzqRk7oN39S2VPUjxDC9G4
Z2Km1R3MXF7KXsui/Hg/4LccSE7+Fzn0XTCYUxrgRXOM0tnTENLQb/ibWtUTngOC72Lltqhs1RqH
z192SXdPyd8v8MljLeeSTEDDbqfGZB9L1AncMd+hV3jWM+zTXKLCsRTvszxNR+SCfjz6p5u7r70e
E+W1rX86HilOhu7genVoesEkIshPHB4aLQy+a9rM0dXZrBpH+5nLF8bFwzgcTbVibB52N3uyJDBT
VvmMJnoMZ3iRIPpt26KTVLdzhKK70dcGte0Ew7LOq3RQzC8s5MOTxLvEcxs0ThPgnTrVdu00+HmU
UzgP7zCCG+n1iCFErURjiUtJhQE0aSUgoUI8wCzqu23DnFyRsm4NGzZWTT06HjmKfAiNo4aNR5eo
nCrsM33Qtl03/skA/o7zzxnNQs5KGQAgDdbX6WejKFfDMtiROL+yQNLMqn1hu0ebn1WSRu7x6THh
ePL1zFA8cFxn9FLQ6BTn6uRovtWshM/9lMIiU/P2O+4wtfYORgjJMd5snHJZDJ44cPEuaVR5mOLe
mxVMXAdkFrUjGIp8pK73auiGbVdXbHxJIhvKZPdXre0IH1jvhdbvNBONoaGHOlZZSQIyMEJGH/ux
755qVq74BlZGqNfOSbE6zpsozirKDm1RY9vRjMiT0XKt8xYcXkoMCE4pgsbLst5IOtTG1xvNxjB/
mrd2ph1UgmLvLWeT52Ny470uBQwYc1Yc0oGJzcVfhvtDUrDNf2MB7/U2/TISC8TDAaUiARfb3oxV
z0lB9h7zTQHJ8YeL8eD5b0iMV27yuTLUxCe9pS23opCArzf+8ybKEa0Ro1IPsxL3+5It3tuX+zz3
XEKkTWtKINw7E3JUc36hsnIcRyXWAJ0bD9vMDVBqWufbR6moktqTeKTKlTjaGad0k7kL8fcpYgxG
e5+NwdMP1ezTK24Z5I8iNXkpIAm2h4ax60c2CePUWBlXsFOOiK//lv76dYb5AmZQyaIqQQsAspOw
Ubtm20cAVrRhCA/GBS2WQixDl1tgEf2/VHzyRO6TTFx1WB12MlHT2ToMMi+slnSNdPNQaz43tRQq
VR1MMIh7YFAY9UIV7pPPY33bVb3y2h5kUmFHFps0tEJUVulEfXtaMK1pY6qAB3MCe+nK4zZ/IfGn
y1bnBmVg+A9AfideILcO2eefVN3W6wYOIorYd5PrURaygPFGAP9B724z7s8wUd2vMWYisqdBPvyj
68Y+4KBJfpn07hDojomuWbOq7+vY7SKXj0JEPdIkNyD+Smyd/wGDiety7V72ksL64oCL4zejF5M4
QCYC17z+EO0IF/4rLxYvxR6iI7szqTVWffe5JsXEeBhOHpHdFwLT1FXwKX2zU8GOC8QOnwxrBTRD
B5lDECK27/KF/yNH8cFmutOpwiR+UJ8sMBgTgamMVh9NoAQc2FoJ+qrtG2sxvPRJmmjGvTXQcQKV
ESlBvAMjQbofoH1wk1e2pQKGujJ6Q4df/gzCfwIOLUVjB4BmHjWeB5ENBcU7x3/1/CAc7/mhq5cz
Jb2ayzDOFF8o7/WX4C/ITXTBXP40DDJFfYwY0oEaqtvyE08nlbtTi7McJJHEvaJWsX37Ewu/jSEM
mftqBfwSdG2/Yxm6Cn7SPKD4fvtPBcUkaNJtfODYyh8Xw44xSf1D+hwcO7b2p9Bh1aJFZ1sczpAq
DpRIdL/iHl/9iPGpyLMXkzjt803B5dYTyQzlLn3J92ocf0JA+BpoNTInbL93TsmFi/dnVeZ3Zwaa
rVMLoc3Lk24o6FUnKMgu7QJfGKCryeEJDY78r3wGoR+6cjPNg3c2TPFiJI1eqDeATRFBmHAhsmqR
ipq6HXvqSOO0B4LvnVfHdDVp/NVlt1wLPhA8xY+BwanTBZtL2bHtWBpQ0mMOZTLjocdHPqxJC8ig
oMa/lUEEwiukPS2lv1Ia2ilhQi/GwaavFeKsBMFzOT4q6Iv8GIL5KWFhdIEM2fSjrxlXRGGjNnfu
UIErz+p59zU4BtEcB+uLmqP6J4bZi4TODBDj2UXP2xRnKRSmqg7kzyi3ThkPI5+3p3h6DUU7MgdJ
czzLHP2n7cA5Hko/KTDRza/4Uf72NFd9tCT6vJNyN1FPPMUowSzIZy0ZZxD2KU47OKlqOuQRaJal
JI26aESz6v7xsTO8l6U9khh9ozS2XN8JwI21GZ0UZ61jEkRyD9baHfDmpTxaM9Gou3ISgXQnwWpA
5PmgXCcIUezRPYCIb0H43w3ybO+K850ANSk42cR46yfTmzGjD8B8eeP46Dxjg888BW+3mNsOo4/y
OskR2u8qIY+Q5dkyb7pYBffPoUP8SMdHrwzo6fu81rdgAyJKn5oyaL5bqahj+8mnOS5YrZqg3zbx
kWpqMmlfHmH5Bm4kOqeQcE4IAEJIEjYFgUsZE8Dgpub8yCBWnxAI5PoXvtaWjGekcyWq3jIR3yhc
DVYxtDPQqtNyBj6LCF3dnMrQyWvTkBSVLemtEhgvP2kuiEEmon1usti9CYaEl/F1BHHMYHKOCSQ4
UkpmyVme/gGZjEOaqIpTK/IkaWlfgwNhpkmwvMCPV/MQ+EJX0DBxJ1o969wMI7jl+UH9+0EcUuRe
Aq7TLqAY1bt6pnpB++6RnKs+txjLUd9/vSqYQyhJcy+QSUdaRw/iHMwlkwD8g7zzwaiQQqTmZlTC
L2W1hA6TdpYQn2krXLQDOEzzPvwXwthS5lzkqSfdGGlNyW85pQ23/wMs9NW09i6OxU4inNIV/Qlx
z02UE/4tMWlytYEILpYRnmpLA/97IISy9M7kgkZtlP1wmQInEVgfAI3tMAENF30KNsWkJdbzHgC1
OVvlckwzld0EoiznZJlpRzN2ddhy5OOv7V4zFqMyNhMC0iLgv34uoYJoixBIWC58HI5wEx/cq3j9
me/hLRZRq6tNqTIb9Wv5Q5ZdGsSOmKLDNklJZfKFZ7XQx2gE54rBsKP60bH8VR7DmTM0LG50tbH4
Px/or89t6wqBBdktcC5wreNT/3DpKVQOcoFjyVmEq0My4MApLYMmZz72ICaiS4tHHRw1vzfV7Nyi
CGp8Sg0vnNN3FOkg3tlv0oLxZiimQ56L1GJFLeVDswjkvESaWy6qHq3fLvH+Fgmk33HJrLyTCYl0
DJ4NSR3OhUisGKalp8XaK3tNpF37sCGJt7012ksbKZvcztczyRW7H0PS0idOUqjTsSVk7cbdiUBo
6dYCZVqoDcf5Ofh/m297ZtnpaF+4Fu9AaX1RbAJ8cdrfsB0kFq/Hi3XxL+CdlDvpcUPA3XaiDdgU
XOCRndy3KkdlYVCs4xrjxSX61dXCFAvjiBs2j1X4wBk9gXj21SxI5lnRSzZmMQj13zxoTsVHj3VM
V2fWqf6aJvx07SSjTE5R38qhScsEAMUvjot3bGJedf8eicC9QHwxkfSbs/qZlKX8+mRfWDmZO1UE
Dekyt+qyMkN2RXgfdH7P1ap3O5Z8nkYs3lbTdqxL0Ou+G04eVR9+5Kp7qiKqes0rSDvTev3P07Nq
m5H5ivebArdngNtkJufXeur+ZwouTwuAlePUOD6XfRNREeqyNAF+bksj9WX0o3lCC5h8Ll3SfpRJ
wUS+oMZD8TF3sobnwKhTxmkMH+MxTxWZvRJ2WhTXOZBPE6CQwiJdxsheK/YoqaQAC6Pzb8yAE3sY
jYMKSoNh5zaIFr0Xi9fxTcpOWtvuxd1UtzEW2HV04+hoKdLL7es8j34T9rKX7Yj+qb4yStiYzWmr
MOdoy3rZVuEZqnff+N1L8eAl980341b69bVvGMCcS0/pNdCZzlLfLohwzI0AH3cZ1TWEOdfgxGJx
Aqwa16EwvdXiNGQe0CuIKcQlYOeb1QLUZ8y+CJBi6Z6p29c5b6lxWwwCjBm/8rT+la5oXvd0eyg5
7HpRszeOMCb8LpVd72OivEY+m/GtY/o/OQYOb80HWbY1eXNSW89VGCshyHw5+DJ4WxkJUcA8NmWg
RfQ5+Vu9P1/Y+3un/xi4OPxuDQeiymNQ6Vkv+RK3SX4ADnt9HCkPXHDP+XawD8Fs9cNeN5TRJ8vl
aqbZZdiysbflxom/kDOhRd612XYxXFS6XXeMZEY3patKUnAwklMOwY5wTR0kXNtEp8sMtVLXhjcH
j8YqaXQgEnLaU0z8FPQNbwCB8iofzQM6QFA6UF5HK4JvstiAxsrANjGEd3KOkbhmmhcR8KC6s18i
yJFe8WG2E6Gfhi4EyWyKbtnauOZIwBhW4Jp90+ug21CA1RJ9xLSZAlrJLHVpyIR0pqXh4GIrT4QK
YuEVRXSfALVKeVekQJFvNp+tfQyumlVbtQapCZggkpAkZ5dk325Vy1LwzxHSACHVGfDju6xyw9gQ
8d6EjNdUn+xHtKcCJREk3LRsxEGIKqBhUUObCgFl/npLc6tzeExw4Lwr/G1TrEXITorKTDU/24TZ
MlxyBdqO1/OwPHRvS3ZSwPonA4nYipQP2aOW1cMoRtCyjQq0PLbAAehX3/vxpxOx82L5zD406MUW
VyQA62gkihovZs+Sux5iMPG1w7ARe0Ok23bYTEcqK3i84NNECjb7W0aj/OyjNBR252DVzzdtYZt9
fZk751X7PmdWgD6q+wOZzQeA9aGbVWm9CLQ8zKNOLuVRY4BqZY48TgTC+MLWG2YbwHX3DDEi4xwS
rsS+PFj3F4jqfJRyUCwUxgQNQ1fjkRELIhNz0zp0olQRYzZeJOdNsc9JSvsdOmpH7uwpNAclMlT9
Nlw6nRat/ZqlWMqyNuvGUyB+KsKW5gwSbcda5ywcnyeSXdKU2THebU9D/oaX/NkDcnxMN6Woq7/M
Ge7eAUz/oYrinGEOa47qEH5SXDavb+r6VMl6vJS7VatPTWVS0a0z3V37/wEC3FDvkLy6qMlT2NWo
gkv56rKLXm22f0KAXWODv6jGflnVf70U/mjfKlwcXm/CwQTnIs2srRiWznYCbgI/3hjquAiy/wB3
0yyz/DmBeQz3/KFA6oXPI5BzqZW0gqIsGBYB43J9QC/5Rm2jdtyYXuRnFbIaC6dx+mDmcLZV+Nnc
E+zllq4ctHKCFnmnzo+HBdaqRRuIsuF9wkXXKuAJPFSAkvyqVvK2hh7oKg/+PpncG3spNoeBEJVo
JhoL0cawx3VwBeYdLh1PUhSVlA2f8gjLxlp+AwUjtcWIFy1dx3SDgSmE4dfdd+iANURo5heSibwH
QAipUKLVESV5W6nXMfWK1rZxy3yE/lmlcBhImbrR3bTykHMfUH1N00ZT9opn09RJd0R6lH1SsLrX
cFICNTpZJJQ3M6oLCoV4GbkTc+PWbpO0rGiSsyQAAnakD5jmdb8nGe/JUYH9CheAGbJ4Xhti7Nn7
CGrAPtpe8r+ZjV0ydjg+AwjHwKyf25UoV+51TOhZVno0Qms7wGX2cpzc9Z/fX9srCrX9yxQ5U9QX
nfaGPayJ52UB1iK9yf/J1eYp4yCINEJ09BhvF8Y5dn5gxI63RyORJI1UznMzWoyLh9npM4LlLiaa
1ddN48Jm+jPYRRFVdCLF/55LLNGPEnKY1hTXhnRSJMe/IKx/spVeB2uLVwDVJ+QFRy44sMsbnL46
FKaWvhVb5JzpbHUqsDHRcIQYltKgpJos9KNlCzdy7mG0TqN91NAdDM03JV/vwMFu3dgmjr4pqTbm
NMJli8t7hV048Ox3LUb5g2YmVjpz7/yYaXxeeNFklzjR2bYsdY5SNOgQXPtMxr1R642DuQeMQiC7
nc/njXGJGF3XbwsanfJnK4snFtLCkm0kEDHGtX8z2iCHUFQlsT8oti3SRyKawAibfr+lusbGh/bm
IPSyImDMS4V1gZGslvRw19K/cHp5fWHB15KyRVIju06dp5caWFx1RvmD5HxIrVx6x/zxuVeI62GG
TBNIpoI3W7DQitZyVVhr8BQcK4R1G7cg4j40UKDXCmS7H4Z78tK8BtTaD4gUYiyWWhv+Q9VqaiBa
AmN4sBnFZFxXabyTLGnPWH1c5JT4C1iZj1ng71sShwXc81z4lpruHm0JzbO3PppLllaK6EvLkK07
VnElePrZTLonX2rhytkGktY/sEfGToA2DHrL38UamQSqqyhQRvS9OVMItZuAB/ejm57spgajWJcO
r0J8/tOY/TxNNx3ddKN6qcLoH1r4ZiEtG5SjtkpHnnvAGVDmbJ2raZH0EQ1i8//lofdvEc3OU6uh
b0HU2P7tzNOiisW1MJ/5jwcs2eoIvRN4Epn8Rz81pQE5YdN4DkCobLV1WWTgi+ZkqbLC6C6kvo0J
3GbWUamk5R82IpddOknReFhkNKE/syXNztKEDYFE5RTI7TNlcONM+/ewmcsTJLn6TuE4MFlnlqA1
gW3UbhLBxwnbwfJsi7J+1YrBJHYOhIOaByqtmKoObIiMUi49P3eGqUPPIX4igLnAgqArEElTibzV
Qt29NNQ2/EAFVtaf5ZsiSq779HvqJ2e7zEHsq47y8Iq+7kHS0Y1Ed3VAfjC16xNpvzBeIAW5eRXS
ohVu910SzKd5VnCAA/Xy9fT/A/7KLmaERgM5xPZnOfQAj3mPEFSdc33QuZeJcdXBI7PUDg2AjDHc
/YJre+iaBMzM165go6i9WMeeIxMhybFUiVUeQk1pSv59ujV77B+GkfqF0Eyd/eeO9UEwiCwCuGhg
37hLcveNoCPEowZHnZXDHjml6EE1x52GDqjxqH5y4q6Ly19PiYIfaJFkrUEYqki4Jtlq8ztwRWRn
Nc7IfASaywfbmI8ovs7+DTALBDue5kmLU9mRj7GXTOyQTrmoihH3HebDQx7w0c3nUM3p1Cds4ugL
vNfVqciZEepRgikVBVYgc8CNBbaaAaMFHHFu3m50ZmTjPC1RRYdWghmjrx6wFj05rJYygh1VwDgM
STxsBLFu+BMj/57R+Td7PjpQSSV8YFAR1tksnzubFLAQum9lHxuewTxJh8iNg7MXugRuG+v5Jbvr
rQtEsdDformt0VeZ6KsvZKqzxyuT67/TXNu3Wow/wP7YszQi4lccZC5npKuyIVHYobRJUfKr3isG
H0oaR76Itt7oytu6fzqcLPtK8CByJ/wMDjHm6OLBEPzVCBLh8vmsfCsEJw1e30P3mr75PfW9wrYW
YRFujVk1HFQ+Xg/wl6YxfVZZ1OULtK29p34sSUrP5W0ro4hBApLqvDyQO0N1G3g2pqp/ixlmT8J7
oFknfZnJE/sD4+tzVS8Xep1ocHJ5o3VpGFOuzHzSjDjtM5lVVMBdf0JzX35oWi2P3a0W6Am/INdr
+2QGONlqNdSmQ8c2TvY6cVkME8MgU9MaF+mo49Z5oHrxi1RSwzp3qxHHRK0Xu7hxh9G1mX6C72mc
D5FhoGhZ7OWaX6xPNryjzcFMdhAACsBLc4kW8DpFm9WxI7ZDnttFXncLOOAto13dOCvdpGNqdVdA
cvPlX6uSKFXAEzyMcSuj76GgCiCjS1LNgfb8E92cPCxyskQaG7yLmGc+CJa4CR/vmzbTKk8q/I/P
4r+5HEpt6qb/viWXl6oUyp1D5E5bm6bc/6gJ2vTSvLPlYOAra7XiZH3WwJ1aHeY+ozARmib9fTst
AK4BpWslyOgzBqyMONzf8sGWqOWA0ZBbSJlIJtg/9sZD/4qAoDCCTrlGyxMAzsmcE6WoRKRbBRYJ
wuso0QrOv914lUbiHRXwCONr7o46lswkKZREBtzH/02gNI95c+sSgER7SyBsXy4h6gte3UVxWa+6
cIOrQYvSuUCOzQchZ3fs5zqMJ+hWHHGSdDp4Fxp21nj3sWwSozOx0uNE9AM3Oprk+RsgixUf23eA
1HUsmLuu2oxFs/V8OJdP/GP+PzoWNa27yd0tPx09uefH5gM8zYIkYmkFwZLmCqfqVLKsgXO8ZcMq
nR71+rOich1ZerRURf5DbMZaX7e2lyBa4ESlTL8Cs/fi1/REeNDVVFxTWujXo9uD4n/zSHKbFlHR
78DJXkCxrXxCgbh/+OXS6unutXhQMn0BuGmmmBxqwf2+lzIiopvmDsK9vhW+cpeu9XlYqhDxUqxw
qzEybw7KK+QMGCgDnYgDiADUAIeiRXkHIB0Ey/wirfHSrupaAO9MmburCaS8V4mLY8vnJiA0IPpM
GgJdeAg12qYu3CXKrndHZLZnt8tFqPLteX962XEYM+MDyq+D6d4PXKu8ByQWVSAoEDA5UKsPkGCq
T1kTxjJIrLfkU0KJq+MCtZyEfzund3ruK7Uwgd58nwEl/8EhTpA4jv8PEtMjganwnDLZsknKYQHo
RHcGQpjeEM9yPHBrj0NFAGEROFFCURBxPmQTatCDGcgRP7xJRFfCUYyZ2DwiRwOZdHZj0YFBTlO/
vDFqkJ0swuHZ1p8LDspMPApfIShfKs7lsIYOK0s4TcoSSLsVH8CucVnUn4svFLji0zvF8cdI3BjP
EiEqC2m8IH52ymceRHaPfmCImfzSpfm8CTW5489qLRQPdHqs4/1YYSvox8UL4StDrdgMU7RMif6j
U/nQJe85+5SgSpl8wG0vQKb2Jw7u+3MAvuqrGU4GMosS5QkE451L/ORjmy4pl71SFvJe8DB0s6F8
kMvPmpO6HtBWTVSvj5kMB3h1jfoyzF7qQCr/lDorgq3fVAxoGjzyO/JdD14MS5G/5UyH15cR36Ba
lzDQ3vZGNVACu2puV679q+220296A4iZPdWtuxEopDeKL7g02asRQsJEupbw5VuNten1996HBVot
gVavKV9Nc+iKcxQdfoUfkW1vwTYzToNyMOQqPBl8KJK8Zv9yBbnZzPGLwQ2VeJwsuyjG9VOnuKGz
k+a9DzYQMpt49r2mjkbkNcJ45GQIV2Ow99fxueTU/C36viS2n9w75YU7t//8P0mJSMS4KlvcdJGm
FqBcZCHFiJ+n1q4f+HbJQATAgjF3GSDx7aIH7zOL+TP5P8mJs+7WfCviEjR7pNSlNskU6II4C8Ia
3S8C1eIpN7V/dkETdJuXBjeb5QPfmEETgwwPyKBlCimalsZXkFctfUyCh+xnWjB1FKTCTV2OB6pN
LaOvT7Y5Oinzz31UH+EXvB/AGhzQTpTm4BnVUjmAtJrSs9nKW2VxKk1bbVIZ/HITl/7OKy2JqfDM
blSRcS0BWUkpSnfupK2Ag0P+szyy+4/97Wp0iE3zu0+cT//THPJ1ftMrPYoPYuSR/sfrAJJ8POSH
TZbXE+2p5h+oAImldi+aJV45XxpToODAyZKuv49VfMoPyvlnACBi7WDErk8EinsquGqf4oDb8weH
Ljbqpz9UYnf6fHAoTY51K577HdfHGCA+eAEoO3CUv1yfXfrMDox2gExUzq4yvvsOh9lRvD3B3AMi
4WGvqbDuQpL1ZFERopuqQTkyYDvy/C5disbO31h3J2vEUo+NgkhYOwT7NaUbmDcAE3fTTKVcYZ4o
PABPIUBXG6jvP52IncGs7XY0TaRPRNZrc1/b1KRU6+KjE3hNW1pzP3EUElYnKIP+tPwjGr5cOeeJ
81UVpPXvIM29jQLMrYpZwy4sWCAHWhrmz34I1Qf1n3nGBrAUTbtV5qIyLwp344H25KsxyTzufoxe
SV3XgCT3qkbJhXin7QS3wtzItxU0qhoHfc4Pkqi/1ERMMI3R+YixnGiY8+5QPgeNBPsORxYmJ63r
aByc669KoBfbBtXY22zSUqZUkKgkpqOwFI4F7mwKr/RnrHPZXUw6nRFulrn0Ilq6x3OIU6LujFtM
WK8CxVRT+8ljWjxuon97hfQGIXGw1+BY5mTIdgpIJdTXsKkWCX8NrQvmF/44q1yc+Nx+bbLSseRE
26qx+iwpKKhIuDfUQ9jg8a05k6TT+jSMajr7niU2fLqbHQJJcIiNZc413v3xOoGwk1zCaElGmoLG
44a64zyaEqH+uEjVaY8NGw14GoKUNaajmynj/ouyX7dnnjKJOxLKzM0KP6G+q06LbwL63whVHJqu
7xjjhx+l4Fj+komZ+NqRfBJY5+QiytFkafVNfnPeHAJ4NynL7xqZlS8Q6rfqw+fBaZxuS+55TKSB
zOh+rL8ivmXa//0kQzFB0kimnxn13ODk8l8QZMLIhT289rJ+FtNcTB4QY5kV93PIcO/u2SkA3Ydt
IIOgxw1pEGXhH1D+bDOEZX6E7ESY3Ocbp+nyqw/TNjAxWXhlpY2pHqu2EPaFBNvnIKDBA6ReD9jT
l+RM3+lw69dpjVhia3I8hux+ZU8SH8SajpUYCCnBRUln/QwvKqPN91owhM07Hl9npqLqfU5DbGvN
C8Fgoe9nXtbPb6r/fzJ1bzOWOLGyJLm0LVfMu0bVvIlkFf1Exp3Vhl5Qm4PdjW5a0W2gRV+MB4ns
pfavQO2WNo+G1KeckoFz8tr/cb5DcZN7nvNd5xe3VXE5jNtdk+SW2Is5Qctqzg5Ka1MuJnQMERpa
lGcYP1wWAvlFnABj+GTHtFUfR5QsFvhqTPePrPWUQz+WyXyjP663pitdBIGKiTgJq+OIUmULHPKw
BNNuvxUz9ZKn8Gb1/7N4rKcfqC1p3fn/TY6cfF3zKQU/9UL85skT17K9thG0GOmb+K6fp6khW1+4
yW8YXG8DWYr8XaToOAcsp7esHx9uxNhI2Fu7jIZ7cARI1YwDTGjm5ZQoaAdPlD3GB8BBv253jDUv
ygl/cjpMwbGdPupKba6/5mwoDpVQ8NnqdnA4uoRAPugl0Fy2oePPb3Q6Fcjj0EKwpa7JUYe/Em4A
36tw93U+0vNcdjbInrtkVRH7FOcskERnaBwbveN1gfo2gnUafbsZi+lyOi2Jaf4F7h6GTUm5f6UP
tQIPlBbo+iMi3dKCQ2+Qk2TmWjq9IqdEzg0uLrCQtnmojxP7aZqoEI5thyvsaWQ2uvcznAgBPoyY
eOBsyF4j/g3Yo/o+xZS8dJ/a2vUxPNrbFKpIuDmhyQJc5YH4UOPT7TJ0CpESF3x2+ptF5VyfSgbs
Nfwugnzo2U9bNE/U7PF/6964G5rgQQG+6p0KXY+gwbaMpy+zRgVWah9kLjWw+Jo1BhdqrrO17Bcu
1jK2CFNWKK6dfUghM9Gqxueb12KoP0GtGlCqHpXfystW25OTfXZDt7NBHb+j+Tdrp7DVRSZuBOwL
OyMo+0sthOxeUSMc2wqw/5zE9MaGxD8Ehba1LyHyp8J+Dv+02Y7BoWja6HkUSLLTD5Pws9KWLVik
vDTIf3XXwdGJH+F5uOESdzZiLFWA+KZlnocN9v05sEwzb7FGfU9p1tQ6YylbTWf5MWJnAqSyj3Qd
fhZNBFYD0sVnlF4QDsbnbYcr/MGrVQ7CDAU13ghIfYdAF4RJzArdv4Uk8dx65x2SXFaWCJWiBmbI
XKBYrRPk5Zcs2izgSFX9pleXyLseMC640aXN3MGK/h9xdxMBqii6qBb2LLaiDqlg4d+8eL8KW3Lw
4LCkfzXEEk3DOFMXniYZcuDxZEXyoXRIr4TwQXpbiHYWB1VKx+KZkpctkCGe92RHaSQ6usEm+27F
dQ4TSZmA4Ps8gRmdabeBdBYycw41dbItuBNxUZxdnzt2D1EABdhJAtfWUJPYcSWVBekQ7urgQ7EA
EcNkQ8r2maf+XnIg0sEpyr/jMaLdFKhtiluaVVcOxZBIWkGk1ocdWYqw6TS05AXI9zq2kvkyIk3c
GmxMMU5GtFqnWww7eJVbifDeRCuF7QpIh4tu8/WTYjj7Rxht1pfE4s0HAmj72eTJJ6JL8SFm0/lT
8tNGoRLMagg1w+V4T9kcjCl0y81w12+8kt3qulB1auS3SUwblBf5pNcYOC16ztFB8p/96RpNqPng
FF/aNdSMHh7CIKSmCWS39jtMGEkoucThcAZbAWa+40jFYcBVZufhl78iJZek7wTevMB3n/lapGoV
kCV55R9gI0qegQlQJv87/KS4UfuZNci1EgfIdiMtE0EdzeTUSTo9rWoHafEfkg1NQEd/f6VzK/V8
4Spqn2RGZfaywvRJCw2mDEfVLNZRj931m0Tjo6p7rUfVrDEvlbnf9R/nQQ2b5lKLBswAc3d9/OZC
JvjyBVfd1J8oNjXipkrJuaZ1U5wG0ybDjwHt7kljNxTfi1WviSh/oDr+J7ZhnI1ywT3JSpu3YddV
A0DEDbN4FGaYcCe70j7QKjeqCW2Wk7TkDdn2MDqlw3LDfTZPc/FC5GLlDvyQRHvZwnvUFvBqf5Ow
sw6NCmuyOpLAQIR8ADh3nCeARQttrFfQbDOarihyrEpOq4lsg1P1zmbs/m0lN5zIegLlLPWjOFH8
yfkemkyDwBAu6Pq6Pw34TmbEUMn//9YNTxuf+E17z3ab7yvJ0hYCcEJ67UTqgR7vv5wUBpFGVs4c
oi2nh4c290PhWB3oMW/HMBhHdBlYvSmg5H7Frmh0rgtP5NPIeuwEMlKRYlrLgVnpq/rBlPN/KTxU
7xjn+Ey3VIWaa3Mb9keFUmIBZzNN1ANNL2zpCyte1EQpPVUQ3tcYJgBFmHvhRAipJ6ZYjb9ieOIO
qyj92LF2JX5Kg6pBpCjeStL5rTDafHohC/KsB5fyD/X2kno88VyCviauC9JzhgdxXyM+YjnApr9m
obCGnZ1/fseXBKLAsupdX7PQMQYSVmY5dIaaarZN3APJB8WwfL7eqmynQvJqarha7j5JP6Z3YBfM
dHqMNnej1CCf85Ymg+/Z37XhFHpNsMWsoC1ua4R9Brb37P3xhxv5Cdh5KHiwIIfz7M2H02UT5IPD
Ij+uWjFF7hiCgsyE1Bql3b1xJ3XD5flUWbdV7UbnE0WpHG8H7vrll7aGG6wRkElwzaLDC5ypo1Lh
MT8cUyZFFGAg6xIkWf2JeQ+D/Pm8HC9SqNCeSK3CrG7rxoFTULrPHiAN1APulXO8oFy7zIqdnJ7D
mfMlkM+p+QUm7jiVTXNoPOatpQlFQe79DdPQ5uj4R/C1AZRYSVTxAz3H5x0zyu+S/Bxgh+uYsns2
+oixBts/ligmG2b1GfI+CxuJdftPLaRtXVjQRzETx/4vL6QSsrGB9bIxpnrzx5W8b5hoqpN/c6ts
7oYf/RNhBjs3IShiT+C7bihx4lJrL/PJ2s/AbeFQJgPxH+/ThdxdTBGPHpy0/RDKBXnEJk/GQcFi
AUOkw3JGMFxqWzKuNDwxa+PzDKGesE/8PrzA9zEf+r9AqpBGos1g0Gv3/lyXI5HMMIdsy8+Cuus4
uAuwrCi0tdU+AK33vf2Q2ARRMy0UQiSlkO6TJRWFX9FsNZYFHWWzwr6OLvcvUeAVTw6Iae096Iku
EueZJIZe5Z31I6ZqVOREWnvi/AV7OxvheX47bppqvN5BkEOd44K5gc4pCvVuoWDNiusyjIgKtLzw
wZr8b96xINwqg3srpDrqMyMu/GPlWqzKlpAKo9tXLOMYIPMMbkbOe4dhJ1046nJMzOiuABBrBFN8
o//6X9CDvXQZYEmI5w+7E7yzBFnnE/rzolCyZrOxHKM4paMWg2VW2elQs4m7roM4dmw/GTp5KinR
DUtrShRZgCahqIfXWkXScNho0OLeu9JbUHLxuQbhUKHCweHl3loTC1R7GiSRB1wWxWAKNS0gAQ3K
8ZLKHI0nHgfskMccg4TThUHc4pU9stlT+Lq7ScllUqQD672qLxNP5dPSVFXAFI9igNQA4MD24R/P
V6Rg4Amqad6jsamR8jkyg31R046eTB9u2HP8X5FQkq40Gwn4fcdfNTCGVN6V/3qKyxttv0Vwwvq9
h6+X1EsnUauQYBraufQ3yYXkqvgeW4I9MQtRrRI6A7GqWXhNliKT2GGTdoFNSmqj9SGbk2vTuGEj
KOk2n6wjjZQx2I75Tr2JUzqljvFNcgQexA5t5T5XxymXiHwqRjvfubg1lhWHeHcKq9sk7l4Rzu7n
W8MQRi0cjgtJALNk2b9U7ZR1qjU5lRL4uSDgKGQjpCQTAOJEp5yzF29aS9JOoet3l/SLa2RV/hVD
jCb2yKQ5xPz8H2Jc6RkPocXeNjGMEenXineinknbu+3eF8Ae3nGCKkjcLVjRk75RLpIlmHuHX5Q4
//dQwWFdxH4MM9qI6NbkD4jaoowGrIiCKzkThQ7ABIpYsyqK74wTQhBpx43qVjfIAC+N+caXc5ku
55npnhqnT8xdYNqfWCsUd/+xUJxPDZXmS+SnqXtZJcrHnKagN4DD9F3EF6E0uX2srz7RAMzthBz6
Xk/CPTG1fCrtD0StVwe5hsdfD6tXw7SoN4kE3+m0IXpQ9i4hqQZ87Tz3MmD/J+FCphK9E+warNdR
yWqyL5Pzf1Vd9MQjIEgPrWwcgBZC1+R6zXpLAus8tOLCFQWxBg3xLhSzlJfKSoQ+SuhETwuLG/hA
CWKddvbD6gQE7zI/mRnpIrqW90bSeSxL330vqxzEH+8LNKsDiJ2MbSeHO0RjX1C2q8kSSja0HEYA
CmhEQXEi63hVdU7CujH9Q7moRDVicMrw94eF8sfj77Hc52+vzwLO76Obj4dbaYe2lWEPxWV/OQnJ
xWTOxPbhJeStkhf8SDVqRmN+0woqhtrplW6iNLQSks+HIH3SGZtRqu7cftce5zFods44Ulap1qEK
RJZrR4SRF8u0RctahF77t4JW9fuv1lYbt5JFKp4OTYPn1K1ElZDDwHybgMkO30yYVyKITugXi7Wd
IMMhhwkCEpYxpyBfoij5O3EA8hm/iCXwUjBF416av+0Qb1BZr3h8eSTs/IFoT94GZPrdX/Vy3r18
oQRKbkYa4y2SNeYJ1yjS5tljCyStoKPhW/70CjFaELRlfPSFuDZSk/kMy76KrVXyrAViNBHlXBFH
uw8MAtMP9q4ExcsWfQjRJv5K9eIElz/QXEjwt8dbrEvExgfYm+oOMDWZNdW4fpxl/d+2FoRWDp4F
Nyxcd/SDu5U2UmuiignIrVyfhoh9g6KBwkHbyVUWpIua9Xo6ILZf/SCM6ivmTq5EDMZ/oBwKL58W
wJek6sMwPCNivJwC5LCgj4jt85FZY+Q8X+vN3FqWvdDarD++A/JLZgb+2+e7x5IJVePpU/Voqcpw
b+7cGpkaeWvKLxQ2wZHwk4Gn43dNFJO9IwAS9Rq0nFDzoyM/zDDP6pm3fxmx1JHUNs9dBnxFYIrv
L+bBrlLr1wKaoe/7X6Ose1+/4zcKGiDPwYDYBN9K88C1Qp0QAkFFrr6fBRensjPgB0WmICM2sAMM
FkDSo8o1TMbQNuB/efvDc9b3sIwcUgnljml5J+6zRdtbeK0cbpyGP5isCrA1LqxywXBO1pSHceZ2
Xx1CVAVeuKgqqRsOqpbOMwjlNj79KDBNvdu6rh81sXMrlqH4Cxp8cOzZHSnWMXjslEyhpiorkpZ/
mbluszhhq0Fk7QwOVqBWXpgnPmc2k5fb84s7hKBKGgSeCnZFkX7yU7TAVrTU1uLBb83mduFmigMB
sr37ogZeWAul+NThJlziH7wNEqFa4rPv7tb9sMDFe+fFEH5gWz2EWYGnW9iqui0Pc38wuZB97cBh
MMsQBZj/4LZ6J5Q6OZUhc4qrCwaBnNUtGmsUegn/SVMDYYTadaK7FDq8SFdjOg6dk2xgTgmI3OCv
0+vm8Iwl6q4P/OtO6kfhiAF+5WlLmuttCQp4k8cMDrDLj9V2/0kIX8RMrGE0Tmf2YS6UhVrVTPrB
1Urs9NsboGGtb4C+o2tABRG0V4lQCv7Qf6gUuNvLBfQtRL0is9l7AH2RFjnN18BkykZ73VvoE/Li
a4wrkTEFcVANN/wpo84zryL1ewF1qdirnvtXvln90Mec4Lobw6OAoSQF0E4NXveMTKHyfsst9xWH
V5hYfwKwZg90yrW7ZdALnx+D1eUyRos6SduwW2jlJKOm6afifjqQyywXR+CaOHxjsONjAdmOnqEt
N5BW3HPLAaETnvE7lfli0kRL4uZ502z3U5jatafRAM4UC2DVCsuuOSCHdKx63J5/Qbl0rvjxRbWy
Um/xBjfKbwKH1Y1+5va7aMhaxhq2o6PtYF/Zb9eyRdys1XG+ztlewcd82FyDhPsOY6+ixbFBzDTr
EqxCLbRrVxJAtqcy5iAUPb+BG4ZASucVg9PHo+43tNHoLnzB+qqRV3Iuqze36oGnUwgPUh5bsEkX
GUOrZaA1Q+h8X18Eam6g9x06oSanZnIen8Zdc4V9WLcJElsBYHobUwkZO+MzkLKKspGiCBUrBPDL
WonYgkKdxi4y/wLHglvw1ehsTQfqtpzihDrr1owTeyzAgVkvpPqeGXA8zHHK1oebMZjdeyZJd6Tl
V2VMoP6WsEXFmVY6Y1r4/85sbkhVwJ7hZnAX2L6vhIWyG+y616igW0blsZWY+MAQLmuY/PmA+jUS
r5GtU2eeniCjeJ0Lqx3tI+Ap9O8GX5FhqSjrhikORrzR3XGht2AmMy+u8GCXG2aFMQ61PECJehsX
unGRqcIbvgLfujI/j7NnZEJ4gNIEAXHF/Cdj8H2thXb7heXLmIqWkmiisTW10hJm90CazKXv+Udl
NXpPBVu9eHHZoL9E1QdcfWmzBmJDU6ncUx0jl7ZcCCkLKPeuN6+NC/9vtzatFMoSeNdAzsDpd+Io
NF9xrGOT4hYX24StuVa6sMP1SwzwwVt+Evk9zugvwXo0du8Se0xhr68JfsMhSklmuFOE7Cw39ECZ
SLymrfbaw1EK1Q2FSlL1YDlohRNsr4Ia1F+z6OUAMiAMcTvvSIVdcihx5CaVdj8xHGmoIj22HyNB
K4SNxwdcRyncN6Zu44MkFMuyHLK7d1TwaoLYu2m2hhivd/8tO+8nWSSBMzvjo58qL5r8Zy0wtIOA
aVTOX01E1wPBn20ce2gPm4FHdjefIMRsBJZpJRMAhfWGwIwszZuWBBZMYv8fuLHOc7J/1T6sSqAE
iUSjX+kQGitsfgHnc5VV5WUdj+x1NlRmOQ3QT4yqo6JL+WT5Te/cPHNbcxKn95OZvruy94fcVGfO
izc8GiHGshDQNW71GTq0dEyJ4oMtjnw17oVsoZIb6ymVH5pYX5ReTS8853CuuYKtgZTLiRQgDxiy
VVYeAT6H4mI1Z8qTneGHNZH4mylWCoRslPTAdJdiypmd4Y2q1HWLMMyqEspNP58SsxodLDSTOQgh
0Cg2aQrIdPDjb8hm+ZdVIkhScotmrpubAO5YP/aES7YOQhsoEUIE2N4mqGL57mN0WILkLT8f+cK3
CRZ16I+SCzOg7JuIXzfCwm/mhIixtV6LNN0NzPzbtCdt7lpmc3paOX9YfRZ4zuUq6oJ+LlGv+8+7
gfE9MSlfb+Nj/QN7ELMSXpVpZXiYrqsLOpfv///g4fiGjfg42h8RyRutk+Kkn8DWX5nnQH94fzxq
MzLxQqHacnBaQuniLCfH1FAbOZMAZ9557zva0M0DUu/K9v5zarRqjmFPdUvtta6McOYk8IJu2aFB
9zaNqVLnzywKdfNIVBUAtmx6K0xiy4u2TL7YNkbaRsrtm1hgm5TyTUMaornJ/fJ0RMHWt82ZpRYX
AMfg4uRxPuuYsI5wTi/2583opsWX1iEGhl/m3THYAb4j9R/SRpjew4usmlL6UYL/uSH6UjdxkEAz
x+XrO+0kxCxknkmhTCPctQB9WPMruPlVmPaNw1CXtIGwLZCjDzjko9ge3EpiA76QiM3Y2m8slHvV
K7g+L/0j4KjpKRebrll4hJprFgcodmI7WZPI1Mfrhujd02EUUk8TDBHu8rJrdxWs2tOALGytDP7x
jhshrKd0m+CrLsJkbxFiffljxGkeLuV792gzlH6Pr7VuPxG4e2b8pZgML0BS4RdYYRURBePsrjcC
4MUSu+WO0HM5ecNnzuUUOPsZJYjlpeLlN9qG6HAfbNQvcmcGpPGTp6JsjswGv2POUUpWqQSfu1yk
RAZt/RxYgB1Dl1RWc+3YkTMxYSSAlJ3wkZYzoa4yOuktxJ5vFEFrEdI8/in3MLWG6ro+dX4vPLyt
n94wSmW3pkynXhvkygOReSJYYAcBYhwcfDUXs5RLLDRld8lBz9Jta2X3eA7r2+e8cEFhheLgGjdy
NqnVfTLkbQIaIBAJDgP5CIRkGRQL5Vlg2AEN1e1d51EUEBV+aIqCR0GuXyBZ7XJxbpwh1v5N3y2E
YNj3xYh7rEbkjjycf/cHLfASCS5KEdxQsM7Rbje4rnboOElZ6hqbBDiO4ZqKJJdK8cxkuLJ4sQFs
zFhvurXihdkE/DTPQJrPiphYIGAoS4Jhqti6A2HIbQcZz1xxqY6+Wcv50Ao87mGjE/LiUiwBJx1h
ZAaN1q/vcabNviOUNhRZzRPujb2iFrIeVdl8EKK5WOdrNX7XEB9NApP7ytGVIk/7sOtIcz1ZY6HB
RHiWoK5nVzu1fceXf8kkJIR1EL2u1GSo2aJ+/ghwmOUpZBPjLY9cRb9Fy6VqNBSBBHEbKaGJ1IL6
CRpAIvTzWDAJhDsxgKCXcIUZU/z4HR6/IN732br02MMWtrMPvV04EfvAcd/fraZ208DIgULoG4ZD
QNJIwfG/3D5CAIq2fSj3UHKLOFC1RmtTmC6PVxcVuZoljR2tccW1Zq5rEaelRyQ88RSPrMjrWb/s
UHOmGnkhGHusBRpYNsfWNNGrb2PhuWCvo2p+mC62EbRJaPl3asQVaWve1ZFC0+h/7FzucxA/oPY9
LWR4ZvFvDXXrvcKzplM7Xzm7sHqI58C0XbY75uxsVAUdLx0iC+99YDfxmAY15bLrN4lMrpQ8o57D
f6eskwAbfuqmycmWlEs6vIKp3F0JNz4boTjVAaxwrCkPjPXQ+ub2PMIS8wJ2/H7NayYGbeHwCpbI
/AHI3uM5eDWCujG0TF+GGRgTIBm8qTpi04X7taYJFhMT7OwOcDkzDClEUphLsuz/CDdqNwkPxhOZ
oGXHcSttPgBwZU6r6TC3ItHXQUEf8UcwIKJ0xJHkBJ40g/c5O525WS9S3Z+8sZVqjmuVW97EBtbE
fyESJoCvnmWe5ajzsGg5r8mCIQ73jMZQs5JUjvFiGyVL66quZ+LCEeisT2Z88SxHPQwsETxQtw5I
FGPiQ1NzkMmQFecIvTvbTAP5FjeDU4JTRn5hIios38E9UHcKBNSTKIomLK/oLI9MRTUGWJriMsPs
/oo612cH17Y+G1Pd0b3S9YCbOA2ua/TxbZ3RggCLmHvyQy0dA9IRjCvxcygq5v9w1gYqhOJ7Zm7M
8O4DJ52hN+M3Ltn/5DWtBOl1l+qCGiXELFTtFf4IwTPD3IzHDElZpXpicBllTSQVIsXE6mYHU6bd
Y+RuPEqLL1wyZZsYi0E4pd2cQN8TY1coW1kmG/mKMFKNhtN0oj+vcBldjXGwCJh6cWpmqrHY/VhI
Zwpm432aWkmPFUBsT+WC497Tp946Vl1oRy9alPH9KtC3KU+gNMC81jQEFbdZrFPd90z6/NBqOnKh
ocwoVo9p5bdwI3+qWCmeuW4ao4fXkuYjqapXPnPjIYXqZxdkoK31RDfTZ9jKqVQt2h4nZMEtqUBY
HuSXZ24NszIr4cwpydF8FrOk49/p6e7noZqEMvdCcg/cd8Qf04zBiIaMRYqAcYRl2vHDAr2k4PSS
LyGRU5HJZ7hx3YUnANMpqhMZO4W7H0FAG6t3L8cPUMyf80qfE/ph8WbBCLR6cdXLlW7fGpv3kchR
9XUyqHhaLCUUJbxzAMhgVp1mIurlTmhyvCxAgryZETxsZUYJoMatTQji3InpI+AM1IKfywJ4hl1o
7e7Zm8cDgze4g4NU9vIFTpD65YegM3hIrehthJ+bJ5iYAzgPnmK1W5UpOT9rAjiKzS4UY6PFeAem
ADWNDFgQXAA/wlyQ2gWuZ3amRF0GhCFM/ll4YGYz0bu6AI1fJF3F3JemVcaGk4YN76epYekTclDa
HgbZzL89dG4y1PmxX0afTkYwjr445KQsaBsYVp8s3/Q9/xiXFgs+5gCzcVpdfZwqmdi/eGSnd2jZ
ZTtBQfARMqBrquqXBuQ1VZmIjoKOmTutXWtcCOKKO/KEMCJWq56DrQ0gGf+Me43IMgle61r9AUZN
eNe4zA2XRI0uUEUMRxg+xPsycjl1JHd3eslNIMLIa+/A398c5JQniV0UI8fAtgQHEXEl2gvrzY0g
90gbkMu+qBxXPzfW3X8nPSLYKhFfoPjp7hOioJ4J52s+WvwUqmMgq3hxRrZ3VFimU7bGPTYVgqOX
0JfGWE/glGav0f6pKBxNoDwZlMIBKvRm1Xe7cDazYJ1OnCyR1YwC3VmmWwj4HJRbKmbDIEiFTLkX
P2x3ptihWwTTFcSiDc9Tnowwa40a1XW18Hg5UemREOa0QPyCZAyubf+iedChUqiIdW8XO210C788
ZIyS6ds3nFsBY3LsvFYzHXQo3zr1fc7JrP69Nm0URGIBEpjku0Tq9r9zCTt6KjWjQoAW9jye3x/m
qm2Ok3PnLWsxATwa9xXecJnm+ZefenUgWvx65CW2ryQSrDj+uBuPoWO2YMLG8nslOKaAvWsO7duE
9f0XJcaV/mY4IjGgdPmiO88olbdT1oS47C3YebcNuRYWfkFQM8wb77HjFMunujDhMXjG1RvV4A0F
cPQces7Key4il0qoHfbTPmvOwsueJ4YXAvPWhoJKmoLjiwwchehfh0ma4IfUB5KIMS1hVqYM4SXf
TL2FR2rFiYOZ2YgBd36V5vGa5z+QQsklmx0yC5rND8MTemzNzN8DcPouu45SaJhbOK8cz/XVKmqp
FWSVUvZztOVHl48hUY/JKh+bptPqy/GgNoramdV/fMW9gcmgOV9RxAopImILPsTNHwD5f1vxfy77
PPOkkksYGTkTLmqCiyLpULS5eMemrd1x8tVCk1laulZygGU4UaHSD1K1cggBWW7PGfy4Wg9vPAQk
DmC3A1GUtd4pMdMNqqrbXSXfy4PpkL7s1LUvCaQGJQepj9OmSsfptjVcZSH9eTtvIbVFnjiU5Lwh
yKuj/WvhxWjhDJWS6wWLw+NiSMJnXYH+XcNfhq0UoW4DP9nmw5spj8rXTB14Nl0y1DQoJ27hi526
3W5Jkl5VPUK7B3l76iKtWLDj7ebIFwcPVuk4UpYS6bdYH/whyPcWJSdDcbK2PfWbSSpH7y7kim3G
zj7ONlD3vIsjV+UkzIec6cmNih4eDwXZ4z6QAhd/c19WJe+BkV+lLJkhVGhpkwPoR6Kc11m38fI4
anrd5r26abpstCYXJfrLB4aqjlWifbggLptygbCAZcxwAnK/+1w/bqU2RIc2Xg1Ca8hfT9lQ/6Zb
J+0acOyK/yiy16BoeqHemj9KYb6Zoudqxg17vkBS77WG7JBCb34YvhxtBo+AuetGs82RQSV9B7Bn
MM7bG9LlxJf9H5UaU7WA51Hxi+oYwrEIY9cfW1ZSGpWwLCkbaeS/eJLr4feH3or4WwwM+IgK+SgQ
tdnNAjE6LIMO5wOI8FluHckFM4ZOOkhh1Khh1wG+g4n95MS1Z6paWooRUmOd+WMBFgMewXEJI9Fl
XNP8fEiHi4z3bOvkINc41eAubcXzz24/YCZmy47SV4TB9U+s1hxSjXtmpOZuZ3jbLHWGhxVG9OG8
lHa4+YYmrG7XrnTjIAVO5wNNVnTMuzR3ofCN9b9qlf3UMmZlJq2IGAIoxYEQh/juoFQm0WQW+PeM
rOdnXgqBTJzMZ7CCj6dywiENVTJHISaczxDcj6fAcnZYovR0hRu8aM0nPcwgiKspTQ7+322bfBy/
ZUHYss5gxncJVNCLCqymV5RSR6L0TDlRyd66D7NDjd7G23EsDoARPS0Cea8rQsTXRHzUCCAUmU94
jxiCiWfb4G/ABBDFUNn+QRpsR35zMMEraGhwlITga8nTHJEOGXB63WxSOQmzHkdT6dHfC2MI5N8K
zlFBHRxEOZUqInt8E2dpsQhRjY10D/tjWNMXNYVluyG9sV4INJK1nnPpXApW5bXqbzGua5AvzLNR
CO9XzTNI5oV+2mQXboJrUIIO+vdcQEMABNcmx59vWFAHnyGljz2n8ri4OAsjmHibRj6VrVMtwN+M
XhpjeDZPcDL2YrQaUf9EnlYc69szvDn3MhW0h9+9XehndNqNCsSwgufQBI2sYF7vbwP2uQ1uvh1N
dYqcXQYAOh98+eUiwWNIgfxLDPNM6Apm0tHo2ZVC2HrG3bygHxNW8WavuPn8TyZHs+sC1KDIFA1n
r4SE9K89PZT/T5ODjmTFzjjGzkFdrguvQpW02+OJRtGlcOvxVw42wfaWsO0r8khEMmk0X2KdSpCj
WuAM0o2kJPfJgcFB6DOHFSU5u4sY4CQI7P8i/s7r4husMtbXEWNL2tr5/EyFvfgEk2MXIcsoiE6U
08cD2BKUzSY0K0KQfqKjqcBt2TAuXskGJo+2lr5xA2+7v/9wbPF5TTpwTRbyvmql+8dqbxJfg72g
IMDu9pvuSKBnw9avVYPjxNNrtJb5iuN+dCqaw2tZMhgAThZXNO3EyclJVWdk6K+G/3bUFIIfm39W
oMyTQCQ5cT5SOs6El3rXXCxHatHj+5NVubynppN0iw2PQ7xrjGqmJeIQShi5Y4CqgV86rg0I2O0z
wtakndcaUJY6pieLTX4Le2440lcrNIojSFqy2Grl4vmzS6VOhVcgthaq8a8YusL8trXqp7rmUee3
OBKKzzTJSPX1UBDfbpVLdqNZ0SHWddnHGMSuGisG3pNFeny7f+PKAMQrZ/Of6lw9lW6GLAx5JGQH
0A+QvqAOSRWa9qmtDtsAPnyBLYX1LtQP6q1kA9sv283xEABkCd2GSoks4ouCiAyzhaogJ1/qBb8G
+6CdD+YYP0Y0DOslN3+NNJ8r01Rc8dam8yzXSR6wBjjQwaP+9+/osQgQbFiAe67GE38bIqxb/AN6
LEXWcTbdqiTryx7TIRcOIC+0HKFghYc5zwd3zI4P7LNM1UqvcGr1y9CFGcudKacfSRUW1GDbhash
XvzOh4oWQ99Sn0kHCp8le22FXWznRIpT4CuPBFgJ1HmXXO5uvsl+hkKbR4h8Hs7VdTtwIxJc8ZIH
RjeoCCcjUwDxfJayn9hdjbt6Ok1exZeeuZ0x8uD2Cgsd7j5h2AvbiZc1HEq1F33dZVp0d0Ntjr+o
GsqFXDmIzsQmcLwu3z6wyxv0P5NJDUGS1JGzXCIsFBZAZmnClyG09aKX+GelAmHSiaTHxsvmrl7O
8rtxwTcnOrby/sqvMZZ+HNBbcf5JMxiKHhWG9BDknEas3XJr4Kj8A2Es+PEgygmFi9fvnwzLNpyM
cH2B58qITC8RSES6bLEAdH4zdo/h58TizEFv2re5JvJtAJ89/c7RQVYwwfzBhSQzpR6QNu2pn5Ru
m9oV7HU5f2j5ihoX6chsD8jrlQAQ1XaMc96PxCFOFLhvvgIP2srfeAMw8LxZubXZwht92Xmq2nIG
KfmfrqL0BDhPMXOqooLSWAKF7EPhuUtmsY3roaPd/m5vRHuyMtbcHFs/MqgBvpYNFYgS1dZogfre
odyiYz4g6iKYMWJPafePBOLoPTKsYhMhgXV9KffoG+Y/LhUyAVDM0A3spnRI+sAptTi38hsmVEqM
o/+juXDz5gwe/gQoVA9BsBQ6rrxxI6BoW2Xjh7eXqM3V+T+IDutOct5gJKd8Py9sBL4SFUK/r4K+
eINjKzbzk89yPT7tLeVap24IIaj/ukRVK8bUUqLEPHSJZTnUeKwuNkKsvRP0e2GaazCvcYzdGC7S
0Lb5+bF/yQQtqxLllnc0a0udcWJq6QGOQ1bOAtvXAwJgF8Jg71zXPe96PazcnqFaIpt3uV8KOZ5u
pSbOmYWNvVye8CA9QIPAzaJV6Z+3XJSh75Mf9YA4zGSYik/RPBhLYivVWsV6rJ58qVat6z0MLzaS
F+/Azv5rRJGx2W5Z+W8RFVFnG9/O3QCsUdLynWoTI573iv9DTrgWwF+C65AIeIWXjg1x16CuUI2F
YN6Qoza0G8urU8ZxAYO0X5PwTA8FKd2hrA7JSC9puQhCovG/oTTi8nvPVsfKRycBLgM94TO3oEuL
EZ5TEIuaLArC1zuBR+H0yzTljAHVhH1IJ5FdzVo5pTU3V2NIQ6WPzBqhKCokmPS+daZjFFBz0PAE
WWMQk7p1kbCPzJzbFU10Q53TxI0SVNI3cTnodW851ye0mevXGHLisZE/mSDYscdNnUUPvLFslq8W
WAhoZNWe8RQ2OqGawxEsYuvRrGiDeyWPGOpcEaWAMRHEPVMfBQHajd69zQNj07Xqe32Zb01/CxHR
BS6crDvxsmS/4tca4nQhepil2STRhWr6D2zqLsQtJ2pdqwVkeDcx36D0U4iJ1zakTyAamlCxRTDI
6PmFSXXPz+887lYAp9EKSDEp0GnFKxq2f662AsiXBZioS5Dl770O4rvxANaSis8jcjklR0d4TfXK
F9llkll5KZB29DPPi9Gh2RNUsmzGL9LQyWP/L+UpbojJUlZ8zuyihT0OfsS6B+WURDTcMv7DIFDe
BUcuYrde69qJQ0iUz+4sMetvgypm1z+Q+lm/IH3F4KPAAKXVl5KtUm1DZSMSH863Lx9dTq5DWmTj
7KRz/8r9Ef2s4pAMCELSR/+Xt2ghZY0I+TJ+TjgSr/PpxLlbbw/gO7D8UMRFr78lAWD+vHL/FBsX
y/CfjCBrwuwCcwBpR2PP2AUZQKrvi3j4Z+CQ1WP00/sm+kbZFCaqNmH3c6O0uEHkQoPtFZ+SyEbQ
mooC7K8eafRd0uuLvXF1/FHZUkXK+OX+cCSKZPNkz38gxmhd/FdOHDOohAOz4Bl4TItmzc7Rdl/l
cERQzJDvavu7N4Q8QHSTyqsf4XxN2Gu5Pu2H5yiGZLBPhBMnmcpYV5zm2BbLYEQId4+4v5GfJGE9
oIuBP9qHhncfjV+/h/7g+vj7TXmg/IWJaI3Q8GkTYqz6eWUUQOEHGlcg7UyhwoudIfgdkYFu4i9+
Wy7oitgEWeCFhgqw9tbda8mH6R2jPLJ/hqGq+mq7qKd3fhlF0GJds2WLyBhvpUl8GekUeljJbgS/
xCxiRxBc3MD+IwkcSphQUQyStELVLnc1R+5Qu9d/bO4kXYS+x9WIgx+9pkEsVByFw31SSV4aSmFs
eBICMAXfH/Groykpy4rCG/Q9xRUMCbt2+5waXXeEWGT/k7WX2uzp1IOd+jZNuXgiGojXIn97lDeF
SVyEIBTPF+EdokYYeWyztcFW2Q9X9eHb1l4xrdABGPf8ix9gCnJtXbvAuzgZImn5HkWqp2G+NWfa
eztzhr2N3Pptuo08VXnnR2Ryu34HhpXc/hx1NbDCxKJFfQhiLfqb2OUHRTUSEbKCBdry6912RXle
YvdrFkvIS7Vad+YurSvwvaG1Pqwvyf/vPpF6KyJPVYXE6/D1uNBW1SgJUVyhzKQvwsX4Zfn9RlT5
MpAmnH+JDk+smmjxHPE/vn8NCKfJ7csq8ZB1Ka6rhzhmfiaOfauoUu8C1jMjUCfP2wvuHdm10OzV
23JorZWs8sFdSXE8NKof/0qOndkzL/qfPywQkkTdOyTTkWVJGRCTHMhqc2T2fqh4bX3Mo8MOEtHV
c2dTt02dSVV1kpFKnT1y58yFMs8RBqtyTritk9WNUrnM8BSRK1GJ81onhVHlLnvppepsRdiS1Ol0
ylmtJBXpPpa2yZUgEQ7S/GRJD6gZ/8JKW8WgfemwM3BF9JasiorWqh8twJaLVeKJ873ZtHUwd/q9
cuADoUv7yeu9//r1CXyxoLH1qYsga5wbHDVPIey4rQWO4vVLeOObata3TuwWDPkQedk47iBEytay
7AyXYXLOdM14eotN/v7Lbz740gsplkXimxc440yoIKfo4wb34R3C45tenhz8GhZ7/x86bHJ9kRfN
oWi3sMYJwD7Eydg+ql9E2UVfhNQk4inphPGYg36oRT7Hspp+eeKjvUp1Z3cFl3k8yVceX2yx04Jj
RYJGlitWleEEeuS1nsUOYw9Cjopiz+dNz7y/nKackxKPq7XEs2W6juEzYs8Eyh3uWld9etpfwf+8
iIRffo9vGHO2tuZtvPafkmIg2Z7AjYJ1tAJLKnoPNxfvF0JbT+AlCjDs+FF6MxNua8gWtd7EtxWT
Yv9sXyq8ca/n+Pg+jKaA9zqmmquTZEPB7BVOCRc377fPAtXQFEA/cmN9ciuLgxdMRyG6iHDB0pqZ
nl47FGJNH1y53/ZitpXp+/kwd4BdnT766jqw5WtvwWbsu8xe/qls0N3UPiasP3ENLDdfGO/4NT6i
86ni2mtCCsRIEvspZW8FnVxP8bRAYi1TeDP8FCPp7NXoGdpbKBO+Mf8D9EZMQFEX3wE9RUdm8K1z
CMe4TpTxQ8E4sC3WH1H19Ly3yrdel9lGguxTQTnYLgsTZOhF16TxBWxnSTXdTH9RBs5ZdaK6ME+0
MUI9UZ30mC8PEqbyayMwWwREzcImHkga9dqPJxEHexvgxDQuSlWSkx4W9ayhch0IYPUnxcjiaYu0
PokCHUZ0qFr50nf58eU5swf5U8nYr4Agmhu9B2s8dwaymcLAvGmExhfqG6CNRrCY3VpXI+RrpP1M
Z02eagaAFw44A9JFHvqzx2N5BafozCfN8yCC5Fopy3+cka5x4oaCG2/6V1goxn4AuArjmN2dNCEf
I8X6YjPjtH2GKu5Ip194pAUAUDiV6I+UrAykiQPy84oxb+Un1z5HNMXmA1WtVGPuPy7rV4Zq2RqW
/xUMI/k5eezEZPUM1CmuLzcDzId2pxkIOh0TB9pryy/Wh0ei0sPe8aUTr7E0eKbaDBErWTtRV+7J
MdoUNCVwH8ifLtga8le58HiZLwCgscWdLvjylVB7Q4JiZWfjuryzV1ZUhx4O3dzXHsr7dxM5nyoo
dESWfeVunR9pq6GW5mSk4G7v+2vYFMfW1ubRgwyah4gxi8fl6sDCNds7ny08XazVKhN76lZBhIeP
SsLjzUMUQL5MMx3aYd27Hp2ItUwwd2iiGyiU97eO7N8APfU1c+17Eua2wnR/ghxUxkY1aeugm9k8
c4QQgGm27R4Y6Q91tsVv5hCF4WUPHnebd24ND9bR5DcX8Al9ftP96fjROEqGhibMP46uW9d/4w77
S7UxoCKyrc5Y9CYXHoi6cSGlw5Aw2aw4ru/rfX4jllt0WJV2C3KuY4vDYzfIK53v8/Ng+5uqz5za
qEbQHlUuapYJJLZCOxC8Ji8rGGmeZxXT0LkDHZSEK+yImQhF2x/hm55LnsH901OXNJUG283PqFp1
1qWkOaKTaJ4axmQ0y/IOX+ooFucg0xcgeiDBHb5zoRUcMmFNoChYIJ7xrT8Uvg3lmHoOVa5KzEXv
gLWBcfnZy+1j2uF0WenSTj0QGpHEIw/txp/vwSNXKeyZPaG887WKrWSx13BSqMh+sU/p/3i73x08
hRabPtKe4gP+cG/UE6CjWhTGvqWpQNtp6zQ8rCViioI6YEsywwD6u0V8CX9K6L38zCPOnrBf0IHw
fvayCZX1ly60XfxraFDRe2CaC8qIW6o1jOoz+MdgacR5qixVtbd9NVubV5YyZyq5ucp6JYJMsOtO
VSfRz9UxL0/NmkFAlPMzMzP3MRysu4Eln2L8F71vPn+eEhEEewUejSWXsaHFgp/UduCr+EHxc1Mq
eLZK9DcHPCI08QmtTZSp+FaVDYURKAVsYYhG5O23kLQwJeMnp8x0kUIWyXuDm3PoljbHB2l1XcKh
so51QNsNCtYjT49t4wYYRGyNlUYu5ThKZm+1pjp8diq6rTz8gj0lTkziGXT44jxkhv8n7O8yL1NF
KYfPzdwecBaqKpMv6Px992IRsCU5Ia3bCtDTP+aznuNeg1SB9u0OqjyPDUkPmMGax64qMmZTLxEX
Ru7m6dfHoayB6m5ESaTCMvzdVCHudrPVTb/xpWs1wnVRQNggtTYi4JQeysnn6uMfnWeETmHJD2q2
eUFBIVA6/Yi2MDbpB2M91oVxvMQXCt9Cl/Tmrzg0VjxfeH9mu47Eo3c5w2UDGKPu7ImLc/oeOT6i
JmBjzkD16bLqjha/52coVTG2OcDwEAKBgQBaGCS6YHgUbV5/la/RakwvkjRReJkOAbsjkptsYWyC
OYDtn7Tk0PfqA+CbPLlDvCJsnK/5xKLSJviCHwnNLCHBcxk7yaFAaHyR2suqwyLKNuxM9EjBvGhe
QBkWw6LVBjxkYZ9Qfav+sYb6kx+Jo53a1Eh2CV9ZpJEx8iqCzUH4nIZNshW5S9u4H6e/f/QAqygi
A5+YuDfnQWHwGGaxcBNw3W87lX5hB9vpk+1ddNIi+u4gVFNfuBwJ9AF8gxPyxgGzOyl7WAaG9rnf
GbEPFrtypWbnsg4PSXJBPcCQ9C+iCLT9pTa4CwJM269LMoCzgXzM/IOniR6Eh2zHa4GXFGuiJTxr
AaadFQ3wCbe6CCfhiCFWig44KmF3KqHd4azOiJktUhIY397xpM6yGKrCvxXorHrAq3KSchanlw3t
PE0H1orOMq9wnUCT5YWAXBk3UdhrC3yWbWcS2LCLNIjE87XuIm4/iWCSYGgjqCekLLDgOfFMoiTb
eo228neeHAVuVyq94WU72XGgojKEdxhAkGSgYNZUbyQzenmP3do2j3XAJStw7I3DXb2j7a99yhGd
h51pfbzjOEIGOuOFfdPTSvWANi6wFZMWbvM9FpOd+CzacVJM6uLcazLv/hrIlOvxiqmrw1qVYLnf
r99k9jmQjpthOthN6LSMjSmPjdoy7G0QLe1DAq6UueXKjVAGRdgFFuGV1G4goCwVcznW3vJ7jKGh
aKNDzxDU3E7zUYvW8zFKyfmng0YYgKmfxiglSq8MUfVTbJzXu9L0tsD9Vlg7sQz5+GulZF1LjKIn
ocyM7b3yuwmRjTGz6YtvZ3a3r1lpfjN+oyCaSwFJVdHixgS1i5DIY5CC4j856sWcFpmNMHeaB4IH
/f0PPAEwHGqVCLkzwJFny0k1tEWPHa/LA0plVvjFM/Dj/tLtH7AyntHjRqS7y2U6L4+9Aoe9b9F9
jgGSwYLj0MYwoG5RHSoGVCtzmwlYtHkmsyDEi0L9NO+9KuZqBqdLpmFtWhVf7OD0GxqumtJhmj71
UT/2L+Q0G2KqNj/R7e/AKzNdgRWhx7EwFWpU7Emxa+wEM1oRp41TXJysLbYzPHcAorfPaT2eoksd
R0Z020rrpEUDK+BhGGr2t64y3BQLdAfVsD7m7xuyLgJiBIqpxHeIyAno/2XVNrOqkjNeD2NE8JEy
zk2uNIIP+1MLf1QWD7QdXkR97QtIq86qqklL4Vcaz4WfJfwWAiyzKjZRkcoyhP0CroflN6f+tGoP
W4jc/OUyuYgvUuVf6jhBWH0KOqPyuIpAkhUQtaNQ9DVvABB1XbBVv6gQZWDvhQmJXqfput9HaHKl
tO5WkBEk6kH5cAZb4SMIKaYifMd1NhbwGXSql6lnQxRfvysppPuGV20fM7wzgHIKe1+SiZp/yxJX
tZ7dfeeiCURAThsVFUecgZrXyo3sqvc4uXX/9Q19qWCob9MbgqERs4tXd85PrXQy5evUqbbtHnPd
35CEmWFbGieI2dIMt9pl0gSWAa/9FkRb51knp6SB9wbGgW9NXAOPaTLGm/zbmRxdHtoWalje98CA
cC9SQ/wNX5HYofezZZuqwmuB6Ywvp+7kYBOrPFE/iZjM5NMm2WcNaXEbVvVreNfUOeVeePNtMdNL
WavPc6c8jgcFNE8CnrmizT32QakxLgmHVxBJVFwmZdFXflgPq/enLCn47QMsUOpkBVaVWyhieiTW
qtgebMDD+NkPHPN9rKZOAaPcA/+SjUdBm3QFzNIXdtUCWh++EUbkNhBAC3auBLOYkC2TqLKaY8/Z
MrR2NMWxXkXzHOhdfYOpx0KqZXhi4B7CF7IXWMhof+axypn6KiAm+EDFgEaya4wkT3A55ogKNbOB
HQYqrU9k+htTd+N7qNodx/7/K5Mb5KzGwQaR3DLw/eP/vwnYcUTroHUR+1J5PIik1AFBtTRZ60NM
cUKfY7zOi8acLs3SUrOTGC866TMZ4aygpwEfNqS3zuiY8D17mVWrYCx+89phIs3feQsQFfb080P3
7Qbvjcw79X4ZwKSOePyokRkA+q1IMhEIm5o1JEnaC7D8AFq0713TIqYJZEqJAmqVZsABZ+VaNc2O
yVmuVW75DfE846VSpTuGhWb3GYu7EOLgna/0wpeQXYC4mEQMKuBiNnr0e/E7Khxkj1bF036Ltmkh
ZX2YPjP7MU1C9hvcvCkb88xI3jQbhS8NfzIvXxX8DaUvjW91jtj7JUQqO/R4TIGngp4vCCHlbqwK
bFqW6W0XbWNmzncCPLyZA6vitkPHqnQEaOUCuLAEn5QrQf2g6Ts2bx4RJegqah+iIjiwMKqb5D0j
TpnSJFN/2M/EGIBnVv+f9Tb0quoa/j94hFeYEyLz73m1EOaYJ5CKoSKDKjCTKe8Xcz1DZi84gIu9
7Q6TmiF2sqJdGH97TsOQyoU/K35PPmkZpCIq22u2Dnvv42L5+pyBoHsIirPVZ+AoQ+ZemhPuNN42
zNJJ8E/RjlaXuQ6BqXek2dz0SDNMDB/lHDh7jcbtTF4GU0205EOYQ6xFo2gwK+vEtzvwuuGPepgV
9y1Mg4Xvje3ZxUDImXoLX/UHf9cY2st7EYWAFphG+fv+1fq/8W7lD0gtaZalSA/xiJgDTSzjjX53
qRd45iizcDrbwz1lYx+ajwEEWpE5iG6sUUPZGqfUtehSlcdGVi9ODFiarGLZDgSNs5Bes8AokTec
HMWcKoUvEk3rZrGXA4fkHNeElA2kPqAx69WE9EQR6coUuNQAVM91gHTCjFddgBTYOmliAIINtjOi
GCa94Xs1jqcyJohtULtutQWetgOwKv8VBpVwjlY0Bbndv1ncTwiXcJe8DOsCiGEnAC7zoexqCurt
88pmyGYuAgdfOaxKHzhgg0b0QtpwuXPjgVOM1ATuygsxsVCkVwzogLu+2B0Z953qf4bGFdp3H+KY
mBTXUUFOq+byS8KLHzylcNC7xMo2LgQXLbpMay/067RN9Spijn1k3M1rokD/lz6Eo2DjH4LbU/5d
3HhoC0eyWPk6ckBhP/W+e1dYTlethryOwBGpFJqHAoFYYBJUTP8j9dnpAMeiNxNe1QIrOtLNNeU4
jJsqHeYZoXUPsdueGLitryX2qvS3QthyPz8wK5yzJgqEex6B4vVp84fY7TsIPeU+PstLTGUEkGBV
yO7aEcA/iKjH4s758EF91RViXyLCt5DwHkk7Dif3Jf6/3nfSOmhTseg7LHxOpxnphjoBhHMs5qbf
xS8ENsryNDoWy1FSKx3NCxckUMiRQ7J+o5ZzcaNSl0j/YEaiP9Vx0MTOJwxrwcgbf51Ear2Ell3g
eQalMrneffZ7SId7ga38ad/8vjnuymOldoJr1pBsxsdhvtLmpjL9hSOyOyEZlIX5FbTZ4/twS4hG
cfFj35BxWFy+JqlM5nR/rm7O/X3ITL/6hf9yfbkFCN9ug5ZWzvUrJVguO36dCoQshtg5Pw2f/ZLW
YSO7DkKvIO1lxTfBg+dT8EOjC9R9KLO5Hw5vVnNGPkAqi1mTnRiG9Iwus6iHRdzSEELR1+7I7Qzl
azeKw5OjODhTuoFHGiwfmZFSt0+BfxOMFSO8Pib5bL3hxeWv2ynwy14IOf+ck1KEH0qbVfRwbcu0
KN3Q0Up+UYYrP2sNlZokY7Ve1K1fclgnlS/nzbrp2PhP2CgQjmTeR3IVIDlICtfH708X/tHT0J3t
virjoadYC3uXWQQQZYaSbfa8E4yK0bvVd3jCW3RO/bbEi+6TdZZdNFavZkCWHqRWvaBIx0IwjxFX
M75AA/oMfNGU5ya3FHQq//eQlXaHWHq0ReGIY9IXsLkAC0RnziA9QlQhk14Ku+OL6nwI5rOlh2+W
Tum30VlBRg22eEqruI29XROSAVoa+CGKcqvCoClxaC4QJSYOR6Nu0laLBAzxcYtyGHf1qej1Wn8U
sjbLi8thu+KXtM5Kg4jEqZqfgrSeiSdPMNa9NucILEd8M5x8b5J/Dg8fvNlWZiMFN6O7MBj3EnjE
3lxZI0IUlAEvwDlI02h24z+CyUs0k0BOat3WEj4difh9sRWuYN+P0cgeEPNPD+MjxeP/mGD9TbPV
aoerfd3wkUBIhMFJXYpo/4XkhjtUc4RSt0Oh6ooYM/tcmRAhSAHWTtX9XEDmClm2RoLtuKs7uRoK
UIdm0/+pHQPciWYdd43ZxCW+Czuqfwf1eHGISJmTEF3lVpZ7TemZuHrZ4w++c6pzMn8Y23KG/c7/
4NEKX1BAlBeoqOmiJPlIg9bosOhHWo5HmPRzTcaIZwjG6yLaNvuX3Jdf6b/yZrzSbht6rD2RyObL
+/nCoS2QIlyycfl7I2GMHW7fsbCfL1uqzlcNz+1lyG4leUH1MG3K5ntiI6e50oO3VSE8QYaB5dNA
bkYq7zo842fAF3xEhS7wtrkExHVM/BRlrDrQkmnJIRHLLqe7qJJIuP9HzkYEBWqGGZ0giPkUoqBd
o59M/gqJB9AGlU2In4CBWfVIeCQj7F/ExVKExk7L7QlA/is/7XzTI+YUTDI2UmybkWP7a/sAPirl
spSGG7oJQBMysGw2yFLpmijlJEEDcO9GeLhTck8G3+39IESDcYikqbUBDF7aLzuT27h+dpvJ+QYR
5K3TBO12gQCHAblgh4gSrJfaDeDTMq9Il/3VAr7oOGgzJQxIpkjvWzzIGay0tNkBqoiOHkYUcvcf
5i858rj4+dO8Pr0KmRBSawW+apW8qvZQxYOKLiKJThQraC4dcxOpGBCt8Ot5jw7CSP8CGodLC1Ee
xPD4sv/Ks8B+aD+6EJUZL0Sjc6zC/mxm8RcSQgVvjEex3IQ82OfzV3hrOLyp0ow3gG6bdfcntonC
cV7ktDJCzNCdmpuqY3nAI5XDyT9vVONRCt+b0ESPRLX2JHorwLW2RMmiZE7K7fv5NMk+vKSk1yyy
qFOnIZl9o9kO5BKRs3a2X1tQkFBtxy8Flw+Ue1uT4pY6MKXBC+25btVv75KQvGJyvfr/bc/q3ZdW
ai0qFtkbX+0dzlRxMkrx4+UKnh60otu0R9cADKZjb7/C25V4uEBNTqi53ip2I6/6nYKAy4/W55Dn
9R3OoqUruLF6THRTnEz5qk9R1Jl0QmctCVyfBbcL2/cy5lckWFzaYhH8BNCN1Y2vDthqO2SFRUaC
mlZB6t1aw0TVvnZOMbZhzoKAvDqhkKQVKNU2JRfCKOYE4PyA0MUHOcD/askyawRp4c/Pi6Fce8TC
meiXmUxPX2biMZqLkcsdgXS38lBIwZZGwb5qrLlxWmwRgzKwoZMT5taAIIg/F7pJHHd4dGMJ4oqS
IoIagmysLvROVoj1tAs8p2GoU44xGoXa8OoerPBkyX0+BGbIn9y2HhjvLXDp8sBz21e7l9x4c9ND
8nvxvtZs27YhYpYM6sxCC1H1voGbmz3I4vKcrM0tYhqi0QuxsG7n71crn3r/i1PBfbUm050+GMwA
CV4SIekJoXZCF7OYgF5YhJv6BRqITM/SaUgT2drtXb+4UpceFMsCPvp/Nj6CNOgiRIrP84+RmGai
2OLB1/KAK77S73JedEXyW0aOUr6NmvhrCoYRapXanZ1D8+qjPn9sqIHuWX9RtS/eRocEzgH3HvSt
K47mLjVOgGm0u/PoaFDWFF85Qm8zd77U56npGq5YHnCksMg7nnAsoGOtMF1g/9yIZT4CcfiEjRI6
VtwhAKeC8t3fOXh9JkJRapOna6qDzs5HvOD11fGurbyuVcqFMbmWT4vh/QprjHBZS2z9/gpKjIta
0IGZZW7mxlCFmlgScPN+/fthzwGQaC2EKuwZCp5LyaEdY/Ngjpl2aUXKkl2Ed7XOYl/D/IcN8915
FQ2ZrKb6WpL4FTnllyffSfqmLq23cIke6JJxKC1erKie8kzvK7Wqe0WqvegHEfzoyWcZ80aiyd9l
MQDPMj04vePmJe4bUsQA0wF9RT2RNyq0v4C2nZqBQaVy8CTIcJeWXSpUJKSYYbvJzA1Ej59rHns7
VUvYMTnJNluZX1aISaMXl9Y9xymtLPdOWUMfmPqLsgP8k3pUYqv+IgT2LI4bgTLYaWMPjyngbsjP
9LXe+Nn4smo2WtlXAiSzCjvjrPFT16mKTfbxmtxJt2hYhJ/yH63lvodxpHT94pOmdDyRJS43Xhkw
c9OfVvUQ0x6Ae8ueo5PIFgKruWgDibSiLgpcTnXvYUkXhEJDWNC12Y7jTGzQYfaBntdzHqQAr2iN
8xOAI0pJxiswZHPh3UKH56IUChSyT5mSh48jp2F3nvyDL1tTPo9hchaezc4CZZvop0x3O5+uNsVC
omtTAqW3wnXyOlR8MRRmOuHCgKVqnqukTFMgoT4Rt9LOndawas3zh31GicZUU7o5YlZ9R6Y83xZL
A9WEIEmytM4YWe/xcIkv2F/4RsHFBqohyBbTRJi1Yg31zcwSqcGYWjzN+uq+4eqOmHD4Q2XOLdU5
s3hluQQYSBWIEbtFIqXTU7KUpe/EyxTXA1asIzpguGXUwa0+FttfVODz7bQAneBx45ibfKxISAsm
3wTfA2+CB6yQhTj+QCyTEZ76k7jTcIlI0t433E6utg3MIcrActZdIQ3JxzfqnRDNLt9vQMAe7tn1
wxY5fjSqGPXSX+jemVdhpQbug93WncVGhGT/HKXkIyMToXMMP9ULviwU+1JAg+0zyTbmpIENtNgI
xanfipZ+TLA2uPjWLkJoNbV3j4kYnkX9wSahvwKel0XPAPmabpg7kM8wU90epLLuN5wWTWZ4Cv3R
JYBdktBB3AM55QNazFVLXbW44uyhYNTdzr4C7XVnmskk0ebr0PdHeBYz1QLraF9z6xMY0/SkhXGw
L/UapSzDlZG2GAtMs0J9kYl1oyhQDEtqfybQcNK64hAmWYg/jSZhN+5dnl0o0jvkEg4wdQIhI49t
AU1DjKovvMaC2XynSRynmNRjSxTubvTYabJNsfcIVMcUq6cEk74cIEu+ArnneW9yH2tusjpMsw9k
nBC+jSbiE6A3W1J+Xy843RDWpKUwOKiU++4qE7Y+c2+Oqnusc0OSrVQ4Q8rffVG+LFiXQFHCyQNc
dnaxtTm5xRh1oeMbEfWvHBCGIA1uUENp/aFc0lTmA+015E1ARD5+gt1oBupNVvY4H+TC2W56tI7T
aqvipcPDaAY8Wq70474BClvjG7Zt01vikhk0uv+PnpDxXCJMTC2G245su69Zsg5ItvOvBbp5616H
H1X47Y0txoWqOHf3xVf6LwxJDrlU3SZxnP/Ii0yh/QaLuNYKUwGm3KzyDgfLrDDdxz8g1vkFLeWl
jcCFNaQr8dN3HiQ9nYGkhi5IJBqZGklQZCXVcvUFUZ2eFgb3FNMvG2NUuzLstLq+5teKHn7ERNNH
UPYfA0jy1IZdRSvb8aB8mQMwNdOb3uGeNIGk2caIZCRpJFMQLZIkcGCXWSNdMk11AYQc2wn/52ng
bFZF9PlwDw0BSNih6ai4RxlIngxKTAVtlwdlwIxWVViyVYd1PIMHLPRLLNq/AJk8FeDd01ogxewo
3bs3m7VIaa0ETcRSmxroNQmX1EyQov8c4e6mbX9WwnMxg8cpy2eJrAOF8HOHy93fkVj5esaywq3r
gbmOy0pLJqdNit6OQuhky8OlXxg8TGFUzSwm+iYG45f+iIi0cLPuFLDwXUgSrFEVZjHQBm2Y5IeO
dumExLDKHlFPbmoypEZrWVTTu3gTkleY+hZz95d1U0C3akLEzQuD6e6E9KQDIjBh1ractDYuJJAp
6A2wi6Bti/BhCCUgsnS11FFvGZNj3+L804HtwEd0Gma0uGC43d0Tvtv5K+ji4YkzmS2ql3bBwuvr
hZ1caQjzINasTY+ThTPntMpbj/jUPqB5tKzhGLGH8IuChz6/X7GPs4zavybV7WxNKCjWjwTgSKD1
cz/Fn2InRrYYtQmJeKqiIrTmBK7R3GlypGiH7yek2cioDl+iwCTQMwtJz+Vm4NWi1k7tsT5UtwJZ
iT8OomHUcPcCvcnyP0RO7tqFygoxhp4ByUHTVqRQIB+RV7WlU3tLfiSVQQyMXskJ5vyEAzI4MTpd
xspaSsxwF+A/rGEkyP/NUL5Rb6alsn6hbXDqTgw37/G1FBVbuIPI7ka+y4jfPWSvzud+BcX0lgl1
uCZs1nQPPI90sFtsKYrWMkVRBkvtyz+GPaTxHHvVYOW+f5CBY+3hwRcDZNzooI7zClb66iN4txCv
/AaF3gbq/mnjKu7rwQnxe68uruCl623H+c9R/nhkqeeBNUpXsquQpOhUjG6aTotuVqy4rJsk6FP/
81nncoZJDvFSCn0WyuBOfDzY3zS+COav9g30drmUZwdzGBemQDcu+kkwKTRsoy+YMNJbpz+g/+/T
eHKCaJL/UuwJpzY9S87zwrvntPS3MTw53gQHol/VzdVljMcCcZQlsXW0SS9tkDzUpF00MQPzWf+7
nnJaS3A4ESea3Lt9DZmrwUoMSdQ3BDHftvENFy99CmJnxiVuKNG1wqH74oqDcUu9pOSjSPNf49Hf
jWBjRD06Chm/xlgMdiG91n+Ys9dXakk16YquIxgoyJePwv278KR2HpzuIMiCLMq1qdSkSiESf1dn
9k1YGXZ93qUh04SL5SvSaaXyHYMyx1x7kcyoP2dIFpOZt5dmEsNpsyA6xCidp+Dkx/qjmRlUY4GN
hivyop5OezM7eDlMesv76Wd5F4oVb7OfCySwTc5L1vqZntSiSx1cYwkEMsAt9NaFPoWfyLGhPkDS
c91Y/2lZqNO7eGPyvzkIJr83cLIjsGJrA7/s6mU7IxmHEnxYzh/ldi8jD4vYqz1nUItYURvFxvTT
L/9tuX2DUoS0OUh7ddqND+CS9B6CbYPYFiQKzxqeJKfG6epTaEnUrIWaTuTN56k++Fy70xX0p4I/
U2Um4lBRMchRGcE8sNRbTb5cwv4DDXVIHwCBNxcx1xkeSrwiyg7rX6G6sBrOcbUwOOWQu/TjGr0O
4kIrqKIq2RgeGfxYWZLNrQTneeo553Lu9iY45/m+ctQSx17040RXN+VLtmxPbf1mS3/+ahTGFdUP
fTx2K+TTtpM1HQcLxAkpPVrZcUbzG+O5idhuAzkG17D9x9LTs2WHFEnXc7MZbrz3sabXT4uNJMhJ
hmFuMqkG2PPKSQEHnLk3s6TMBMmTcoklGkLm0InC9PeagVj9q0nYIs72anF5SEYJQaGlAvYw/K88
b5zfeLm16L3KycaJ3j0dheqSO3OhExuZ/GCHjCNamJhvZOGgbrvGaKeCEwPVF6x0CpVaXrRfroAL
D/A6M8MPhSCasgwVLbmZYanLV8oONqNzsVYm9XSwyZO3WSl4Qw2DEJB9ylokrWsJo1Um2LCDBcBw
xV9C0sD2+dmpL5eHcNH2nrgUaYdgP0XEpMFd/ZWq/Pmm8+QNFl9LVOBwr0W52MhhXbEEZlvRAOIi
/gfrexnwi5tVQpjK4WxukkqWgCxSwhKR7+LlBAJQNdrBMbdJHNUDlArtSsvBW9uanN5SBEgQvgfX
J8iSUB4m26BSE6uOMTxbfdRsU11yO10yxcIh5EsgFz804SMygVwv8V7rnWNfUBVwyWCaExw4o25v
+lbxGRX/ljPoNs6ElXZvNeC1YCNE8FVt14lw/9f23Nibhy7uOKYBYAUXf7i7J0S42Y5vneIeFlH9
pASAZnak7wBnwn80vT0Mt4oiaP7gPgMobsXKia1h1GQaqyZs/O7QhHq8H6xcRUjXkgQEmWnyQF7q
N624y5IsZO+p1qWscBvDm/V0EuX0JeZEgpMHMCgFcZUnMBVlphVgJGWt4ihGKE2wL9QEZtv83l3X
ha6R3GMGceIDzd4WtY2dIesNwPF9V7iYSRoEwMyG7XqI8DU5pUuzHxTKX1HYBo0I4WF3Z810dxlr
F0GVX2bmqa6f2hL7AKsOcZrAfK/c87dLqEZu16KlOnISayfRMSX5iagUpoWYxdoNIHNBLJd1OxwX
v9nT7ZJ5dGc6dCC+P0B0C2JGcNUhvDlDl8N+M9t7oPR57Y6t1xGvHRlfLj/x+qonfQCq2P8Crheq
vrB2zAb+Mop/puNwnNfm81x3K6bwBMYCV4VbZQo0q3sVTBGs7NvRs0p1Dzneau3qlb83Uwc+pvuh
FlPpL4WGkUF6cRNiMoOXBZQmxVLE5nTnFM3VIclonzfHmysb15/B3ez4CAbycn+0VbizQSwyvMKg
QyEm5D9RSRZUYHfkCRvxvgfT+E2we+3RCFJBCagwtHzKvB2hkCrL5aHRle0VicsvmfoNBkpBc+Li
4gkplYiXedam6tH2R290t8PKQQNWqaZ5BQRqma+JWU5YgPkroIQnl5TCVGs4cIBtmMEA88LvEQLF
6xR0FwHEK5tsP92RV1dq2bpcOp+KzkE9oEVNXHOuzts/A8Ea2HXSTXsSqocaK0Rz/phoftcYv7NQ
WzvIieqKrLNf8f/60Cy1xWq4hIRSUnqkiu+gxsID2/0Wkfyro4ayktc+NvK6933+Ko60hde8il+y
agFDSuMmzIu4ScZP8rY+O6PZegpQiFR3lDgvA590Pd4jhwy5sp9JzVPDCPpcBl2kAQ2ZgiyX9ia/
+SLse5dMa5wFfWz80+BeRbuvH2+W20InDG+7pdLXAIpwjFr0ty1y4rkwIpLB7lmTp+JQzVjQSGFz
ufskOmHs2Hite7JO3THVLfVs10w95nFgf49nouTONCw8y2AEqwOFlBCnD9+HTiDyGc0MwfDTLdp8
LDkKlRPLIY0yBdm7lzZ+X9wgRB+aVV1+OJ4ML+WqpJ7kOgoFUiq6rrWmy73Ze/hieQ04RyKF84nM
VGE76ozIOTPnBEk8LR+EMeACkZ72op8o9AaI2/61eUYgFZ5h4iE+eWTI/rOTiq+z1HV0nwXUnMSg
x+nv6pgc+dvqtymiA0gCqiDh/y4T6YwVsLMHHmrlKmZpXr7cKiMJxI8fUsu5ZVMiKvHv8U9368//
wW2wp4tpmOnaer2ICgbvwlUZRI5TL8L7f4TZd+jKncbQwJx6Y1acoIrpTI+f7qQ3s7KcpWpfxh/N
TNkliEnCLKk3BrC3ZAOAwBGobixb9MRhIjOtX9lB2OB+Q9PcoNU12rI0aShSJPr6EniWGczg4Nse
39hYg5YXyGTVCWg56eDffL5akbWFSn0tIGAZkpBDzAkg6QrSbsmf8fSO8h1TRIYGPxJML5wqmIyz
rROONssBiFvDrbJjbXuqVUtIUQwuJqiv7AsMPSAxpCtmbUg+/XeRhoeBsQ9U8EmyNApFny4KZPm/
iRQnhgoY3WNBqUs3c0eNHHftjNcuvHsBtJLPcheUbgvZ
`pragma protect end_protected
